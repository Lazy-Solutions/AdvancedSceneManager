{"api/AdvancedSceneManager.Callbacks.ISceneClose.yml":[{"uid":"AdvancedSceneManager.Callbacks.ISceneClose","name":"ISceneClose","href":"~/api/AdvancedSceneManager.Callbacks.ISceneClose.yml","commentId":"T:AdvancedSceneManager.Callbacks.ISceneClose","fullName":"AdvancedSceneManager.Callbacks.ISceneClose","nameWithType":"ISceneClose"},{"uid":"AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose","name":"OnSceneClose()","href":"~/api/AdvancedSceneManager.Callbacks.ISceneClose.yml#AdvancedSceneManager_Callbacks_ISceneClose_OnSceneClose","commentId":"M:AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose","fullName":"AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose()","nameWithType":"ISceneClose.OnSceneClose()"},{"uid":"AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose*","name":"OnSceneClose","href":"~/api/AdvancedSceneManager.Callbacks.ISceneClose.yml#AdvancedSceneManager_Callbacks_ISceneClose_OnSceneClose_","commentId":"Overload:AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.ISceneClose.OnSceneClose","nameWithType":"ISceneClose.OnSceneClose"}],"api/AdvancedSceneManager.Callbacks.ISceneOpen.yml":[{"uid":"AdvancedSceneManager.Callbacks.ISceneOpen","name":"ISceneOpen","href":"~/api/AdvancedSceneManager.Callbacks.ISceneOpen.yml","commentId":"T:AdvancedSceneManager.Callbacks.ISceneOpen","fullName":"AdvancedSceneManager.Callbacks.ISceneOpen","nameWithType":"ISceneOpen"},{"uid":"AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen","name":"OnSceneOpen()","href":"~/api/AdvancedSceneManager.Callbacks.ISceneOpen.yml#AdvancedSceneManager_Callbacks_ISceneOpen_OnSceneOpen","commentId":"M:AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen","fullName":"AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen()","nameWithType":"ISceneOpen.OnSceneOpen()"},{"uid":"AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen*","name":"OnSceneOpen","href":"~/api/AdvancedSceneManager.Callbacks.ISceneOpen.yml#AdvancedSceneManager_Callbacks_ISceneOpen_OnSceneOpen_","commentId":"Overload:AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.ISceneOpen.OnSceneOpen","nameWithType":"ISceneOpen.OnSceneOpen"}],"api/AdvancedSceneManager.Callbacks.SplashScreen.yml":[{"uid":"AdvancedSceneManager.Callbacks.SplashScreen","name":"SplashScreen","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml","commentId":"T:AdvancedSceneManager.Callbacks.SplashScreen","fullName":"AdvancedSceneManager.Callbacks.SplashScreen","nameWithType":"SplashScreen"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen","name":"DisplaySplashScreen()","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_DisplaySplashScreen","commentId":"M:AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen()","nameWithType":"SplashScreen.DisplaySplashScreen()"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Callbacks.SplashScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"SplashScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Callbacks.SplashScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"SplashScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen*","name":"DisplaySplashScreen","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_DisplaySplashScreen_","commentId":"Overload:AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.DisplaySplashScreen","nameWithType":"SplashScreen.DisplaySplashScreen"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Callbacks.SplashScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.OnOpen","nameWithType":"SplashScreen.OnOpen"},{"uid":"AdvancedSceneManager.Callbacks.SplashScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Callbacks.SplashScreen.yml#AdvancedSceneManager_Callbacks_SplashScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Callbacks.SplashScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SplashScreen.OnClose","nameWithType":"SplashScreen.OnClose"}],"api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml":[{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections","name":"OpenStartupCollections","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml","commentId":"T:AdvancedSceneManager.Core.Actions.OpenStartupCollections","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections","nameWithType":"OpenStartupCollections"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress","nameWithType":"OpenStartupCollections.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.#ctor(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"OpenStartupCollections(SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections__ctor_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Actions.OpenStartupCollections.#ctor(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.OpenStartupCollections(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"OpenStartupCollections.OpenStartupCollections(SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning","name":"pointlessCollectionWarning","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_pointlessCollectionWarning","commentId":"P:AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning","nameWithType":"OpenStartupCollections.pointlessCollectionWarning"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"OpenStartupCollections.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.reportsProgress","nameWithType":"OpenStartupCollections.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.#ctor*","name":"OpenStartupCollections","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenStartupCollections.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.OpenStartupCollections","nameWithType":"OpenStartupCollections.OpenStartupCollections"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning*","name":"pointlessCollectionWarning","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_pointlessCollectionWarning_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.pointlessCollectionWarning","nameWithType":"OpenStartupCollections.pointlessCollectionWarning"},{"uid":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.OpenStartupCollections.yml#AdvancedSceneManager_Core_Actions_OpenStartupCollections_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenStartupCollections.DoAction","nameWithType":"OpenStartupCollections.DoAction"}],"api/AdvancedSceneManager.Core.Actions.SceneAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneAction","name":"SceneAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneAction","fullName":"AdvancedSceneManager.Core.Actions.SceneAction","nameWithType":"SceneAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress","nameWithType":"SceneAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.openScene","name":"openScene","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_openScene","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.openScene","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.openScene","nameWithType":"SceneAction.openScene"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.scene","name":"scene","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_scene","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.scene","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.scene","nameWithType":"SceneAction.scene"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.collection","name":"collection","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_collection","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.collection","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.collection","nameWithType":"SceneAction.collection"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.progress","name":"progress","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_progress","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.progress","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.progress","nameWithType":"SceneAction.progress"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.isDone","name":"isDone","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_isDone","commentId":"P:AdvancedSceneManager.Core.Actions.SceneAction.isDone","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.isDone","nameWithType":"SceneAction.isDone"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback(System.Action)","name":"RegisterCallback(Action)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_RegisterCallback_System_Action_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback(System.Action)","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback(System.Action)","nameWithType":"SceneAction.RegisterCallback(Action)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback(System.Action)","name":"UnregisterCallback(Action)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_UnregisterCallback_System_Action_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback(System.Action)","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback(System.Action)","nameWithType":"SceneAction.UnregisterCallback(Action)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback(System.Action{System.Single})","name":"OnProgressCallback(Action<Single>)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_OnProgressCallback_System_Action_System_Single__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback(System.Action{System.Single})","name.vb":"OnProgressCallback(Action(Of Single))","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback(System.Action<System.Single>)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback(System.Action(Of System.Single))","nameWithType":"SceneAction.OnProgressCallback(Action<Single>)","nameWithType.vb":"SceneAction.OnProgressCallback(Action(Of Single))"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgress(System.Single)","name":"OnProgress(Single)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_OnProgress_System_Single_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.OnProgress(System.Single)","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgress(System.Single)","nameWithType":"SceneAction.OnProgress(Single)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.Done","name":"Done()","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_Done","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.Done","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.Done()","nameWithType":"SceneAction.Done()"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.Done(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Done(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_Done_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.Done(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.Done(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"SceneAction.Done(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_ToString","commentId":"M:AdvancedSceneManager.Core.Actions.SceneAction.ToString","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.ToString()","nameWithType":"SceneAction.ToString()"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.reportsProgress","nameWithType":"SceneAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.DoAction","nameWithType":"SceneAction.DoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.openScene*","name":"openScene","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_openScene_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.openScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.openScene","nameWithType":"SceneAction.openScene"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.scene*","name":"scene","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_scene_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.scene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.scene","nameWithType":"SceneAction.scene"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.collection*","name":"collection","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_collection_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.collection","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.collection","nameWithType":"SceneAction.collection"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.progress*","name":"progress","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_progress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.progress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.progress","nameWithType":"SceneAction.progress"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.isDone*","name":"isDone","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_isDone_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.isDone","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.isDone","nameWithType":"SceneAction.isDone"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback*","name":"RegisterCallback","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_RegisterCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.RegisterCallback","nameWithType":"SceneAction.RegisterCallback"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback*","name":"UnregisterCallback","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_UnregisterCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.UnregisterCallback","nameWithType":"SceneAction.UnregisterCallback"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback*","name":"OnProgressCallback","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_OnProgressCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgressCallback","nameWithType":"SceneAction.OnProgressCallback"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgress*","name":"OnProgress","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_OnProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.OnProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.OnProgress","nameWithType":"SceneAction.OnProgress"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.Done*","name":"Done","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_Done_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.Done","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.Done","nameWithType":"SceneAction.Done"},{"uid":"AdvancedSceneManager.Core.Actions.SceneAction.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Core.Actions.SceneAction.yml#AdvancedSceneManager_Core_Actions_SceneAction_ToString_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneAction.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneAction.ToString","nameWithType":"SceneAction.ToString"}],"api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction","name":"SceneLoadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneLoadAction","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction","nameWithType":"SceneLoadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","name":"SceneLoadAction(Scene, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction__ctor_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SceneLoadAction(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneLoadAction.SceneLoadAction(Scene, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction(ByRef System.Boolean)","nameWithType":"SceneLoadAction.BeforeDoAction(out Boolean)","nameWithType.vb":"SceneLoadAction.BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneLoadAction.DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo(AdvancedSceneManager.Core.SceneManagerBase,UnityEngine.AsyncOperation)","name":"GetOpenSceneInfo(SceneManagerBase, AsyncOperation)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_GetOpenSceneInfo_AdvancedSceneManager_Core_SceneManagerBase_UnityEngine_AsyncOperation_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo(AdvancedSceneManager.Core.SceneManagerBase,UnityEngine.AsyncOperation)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo(AdvancedSceneManager.Core.SceneManagerBase, UnityEngine.AsyncOperation)","nameWithType":"SceneLoadAction.GetOpenSceneInfo(SceneManagerBase, AsyncOperation)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","name":"SetPersistentFlag(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_SetPersistentFlag_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"SceneLoadAction.SetPersistentFlag(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Core.SceneManagerBase)","name":"AddScene(OpenSceneInfo, SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_AddScene_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneLoadAction.AddScene(OpenSceneInfo, SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.#ctor*","name":"SceneLoadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SceneLoadAction","nameWithType":"SceneLoadAction.SceneLoadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.BeforeDoAction","nameWithType":"SceneLoadAction.BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.DoNonOverridenAction","nameWithType":"SceneLoadAction.DoNonOverridenAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo*","name":"GetOpenSceneInfo","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_GetOpenSceneInfo_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.GetOpenSceneInfo","nameWithType":"SceneLoadAction.GetOpenSceneInfo"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag*","name":"SetPersistentFlag","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_SetPersistentFlag_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.SetPersistentFlag","nameWithType":"SceneLoadAction.SetPersistentFlag"},{"uid":"AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene*","name":"AddScene","href":"~/api/AdvancedSceneManager.Core.Actions.SceneLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneLoadAction_AddScene_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneLoadAction.AddScene","nameWithType":"SceneLoadAction.AddScene"}],"api/AdvancedSceneManager.Core.Actions.yml":[{"uid":"AdvancedSceneManager.Core.Actions","name":"AdvancedSceneManager.Core.Actions","href":"~/api/AdvancedSceneManager.Core.Actions.yml","commentId":"N:AdvancedSceneManager.Core.Actions","fullName":"AdvancedSceneManager.Core.Actions","nameWithType":"AdvancedSceneManager.Core.Actions"}],"api/AdvancedSceneManager.Core.CollectionManager.yml":[{"uid":"AdvancedSceneManager.Core.CollectionManager","name":"CollectionManager","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml","commentId":"T:AdvancedSceneManager.Core.CollectionManager","fullName":"AdvancedSceneManager.Core.CollectionManager","nameWithType":"CollectionManager"},{"uid":"AdvancedSceneManager.Core.CollectionManager.op_Implicit(AdvancedSceneManager.Core.CollectionManager)~AdvancedSceneManager.Models.SceneCollection","name":"Implicit(CollectionManager to SceneCollection)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_op_Implicit_AdvancedSceneManager_Core_CollectionManager__AdvancedSceneManager_Models_SceneCollection","commentId":"M:AdvancedSceneManager.Core.CollectionManager.op_Implicit(AdvancedSceneManager.Core.CollectionManager)~AdvancedSceneManager.Models.SceneCollection","name.vb":"Widening(CollectionManager to SceneCollection)","fullName":"AdvancedSceneManager.Core.CollectionManager.Implicit(AdvancedSceneManager.Core.CollectionManager to AdvancedSceneManager.Models.SceneCollection)","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.Widening(AdvancedSceneManager.Core.CollectionManager to AdvancedSceneManager.Models.SceneCollection)","nameWithType":"CollectionManager.Implicit(CollectionManager to SceneCollection)","nameWithType.vb":"CollectionManager.Widening(CollectionManager to SceneCollection)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.op_Implicit(AdvancedSceneManager.Core.CollectionManager)~System.Boolean","name":"Implicit(CollectionManager to Boolean)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_op_Implicit_AdvancedSceneManager_Core_CollectionManager__System_Boolean","commentId":"M:AdvancedSceneManager.Core.CollectionManager.op_Implicit(AdvancedSceneManager.Core.CollectionManager)~System.Boolean","name.vb":"Widening(CollectionManager to Boolean)","fullName":"AdvancedSceneManager.Core.CollectionManager.Implicit(AdvancedSceneManager.Core.CollectionManager to System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.Widening(AdvancedSceneManager.Core.CollectionManager to System.Boolean)","nameWithType":"CollectionManager.Implicit(CollectionManager to Boolean)","nameWithType.vb":"CollectionManager.Widening(CollectionManager to Boolean)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.opened","name":"opened","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_opened","commentId":"E:AdvancedSceneManager.Core.CollectionManager.opened","fullName":"AdvancedSceneManager.Core.CollectionManager.opened","nameWithType":"CollectionManager.opened"},{"uid":"AdvancedSceneManager.Core.CollectionManager.closed","name":"closed","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_closed","commentId":"E:AdvancedSceneManager.Core.CollectionManager.closed","fullName":"AdvancedSceneManager.Core.CollectionManager.closed","nameWithType":"CollectionManager.closed"},{"uid":"AdvancedSceneManager.Core.CollectionManager.current","name":"current","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_current","commentId":"P:AdvancedSceneManager.Core.CollectionManager.current","fullName":"AdvancedSceneManager.Core.CollectionManager.current","nameWithType":"CollectionManager.current"},{"uid":"AdvancedSceneManager.Core.CollectionManager.previous","name":"previous","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_previous","commentId":"P:AdvancedSceneManager.Core.CollectionManager.previous","fullName":"AdvancedSceneManager.Core.CollectionManager.previous","nameWithType":"CollectionManager.previous"},{"uid":"AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2","name":"OnAfterDeserialize2()","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_OnAfterDeserialize2","commentId":"M:AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2","fullName":"AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2()","nameWithType":"CollectionManager.OnAfterDeserialize2()"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean)","name":"Open(SceneCollection, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Open_AdvancedSceneManager_Models_SceneCollection_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.SceneCollection, System.Boolean, System.Boolean)","nameWithType":"CollectionManager.Open(SceneCollection, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Reopen(System.Boolean)","name":"Reopen(Boolean)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Reopen_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Reopen(System.Boolean)","fullName":"AdvancedSceneManager.Core.CollectionManager.Reopen(System.Boolean)","nameWithType":"CollectionManager.Reopen(Boolean)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Close","name":"Close()","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Close","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Close","fullName":"AdvancedSceneManager.Core.CollectionManager.Close()","nameWithType":"CollectionManager.Close()"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Toggle(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Boolean})","name":"Toggle(SceneCollection, Nullable<Boolean>)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Toggle_AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Toggle(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Boolean})","name.vb":"Toggle(SceneCollection, Nullable(Of Boolean))","fullName":"AdvancedSceneManager.Core.CollectionManager.Toggle(AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Boolean>)","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.Toggle(AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Boolean))","nameWithType":"CollectionManager.Toggle(SceneCollection, Nullable<Boolean>)","nameWithType.vb":"CollectionManager.Toggle(SceneCollection, Nullable(Of Boolean))"},{"uid":"AdvancedSceneManager.Core.CollectionManager.IsOpen(AdvancedSceneManager.Models.SceneCollection)","name":"IsOpen(SceneCollection)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_IsOpen_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.IsOpen(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.CollectionManager.IsOpen(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"CollectionManager.IsOpen(SceneCollection)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.CanOpen(AdvancedSceneManager.Models.Scene)","name":"CanOpen(Scene)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_CanOpen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.CanOpen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.CollectionManager.CanOpen(AdvancedSceneManager.Models.Scene)","nameWithType":"CollectionManager.CanOpen(Scene)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.Scene)","name":"Open(Scene)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Open_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.CollectionManager.Open(AdvancedSceneManager.Models.Scene)","nameWithType":"CollectionManager.Open(Scene)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.OpenMultiple(AdvancedSceneManager.Models.Scene[])","name":"OpenMultiple(Scene[])","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_OpenMultiple_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Core.CollectionManager.OpenMultiple(AdvancedSceneManager.Models.Scene[])","name.vb":"OpenMultiple(Scene())","fullName":"AdvancedSceneManager.Core.CollectionManager.OpenMultiple(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.OpenMultiple(AdvancedSceneManager.Models.Scene())","nameWithType":"CollectionManager.OpenMultiple(Scene[])","nameWithType.vb":"CollectionManager.OpenMultiple(Scene())"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Close(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Close_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.CollectionManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.CollectionManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"CollectionManager.Close(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.CollectionManager.CloseMultiple(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"CloseMultiple(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_CloseMultiple_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.CollectionManager.CloseMultiple(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"CloseMultiple(OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.CollectionManager.CloseMultiple(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.CloseMultiple(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"CollectionManager.CloseMultiple(OpenSceneInfo[])","nameWithType.vb":"CollectionManager.CloseMultiple(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.CollectionManager.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Core.CollectionManager.Implicit","fullName.vb":"AdvancedSceneManager.Core.CollectionManager.Widening","nameWithType":"CollectionManager.Implicit","nameWithType.vb":"CollectionManager.Widening"},{"uid":"AdvancedSceneManager.Core.CollectionManager.current*","name":"current","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_current_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.current","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.current","nameWithType":"CollectionManager.current"},{"uid":"AdvancedSceneManager.Core.CollectionManager.previous*","name":"previous","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_previous_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.previous","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.previous","nameWithType":"CollectionManager.previous"},{"uid":"AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2*","name":"OnAfterDeserialize2","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_OnAfterDeserialize2_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.OnAfterDeserialize2","nameWithType":"CollectionManager.OnAfterDeserialize2"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Open_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.Open","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.Open","nameWithType":"CollectionManager.Open"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Reopen_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.Reopen","nameWithType":"CollectionManager.Reopen"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Close_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.Close","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.Close","nameWithType":"CollectionManager.Close"},{"uid":"AdvancedSceneManager.Core.CollectionManager.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_Toggle_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.Toggle","nameWithType":"CollectionManager.Toggle"},{"uid":"AdvancedSceneManager.Core.CollectionManager.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_IsOpen_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.IsOpen","nameWithType":"CollectionManager.IsOpen"},{"uid":"AdvancedSceneManager.Core.CollectionManager.CanOpen*","name":"CanOpen","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_CanOpen_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.CanOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.CanOpen","nameWithType":"CollectionManager.CanOpen"},{"uid":"AdvancedSceneManager.Core.CollectionManager.OpenMultiple*","name":"OpenMultiple","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_OpenMultiple_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.OpenMultiple","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.OpenMultiple","nameWithType":"CollectionManager.OpenMultiple"},{"uid":"AdvancedSceneManager.Core.CollectionManager.CloseMultiple*","name":"CloseMultiple","href":"~/api/AdvancedSceneManager.Core.CollectionManager.yml#AdvancedSceneManager_Core_CollectionManager_CloseMultiple_","commentId":"Overload:AdvancedSceneManager.Core.CollectionManager.CloseMultiple","isSpec":"True","fullName":"AdvancedSceneManager.Core.CollectionManager.CloseMultiple","nameWithType":"CollectionManager.CloseMultiple"}],"api/AdvancedSceneManager.Core.Editor.yml":[{"uid":"AdvancedSceneManager.Core.Editor","name":"Editor","href":"~/api/AdvancedSceneManager.Core.Editor.yml","commentId":"T:AdvancedSceneManager.Core.Editor","fullName":"AdvancedSceneManager.Core.Editor","nameWithType":"Editor"},{"uid":"AdvancedSceneManager.Core.Editor.scenesUpdated","name":"scenesUpdated","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_scenesUpdated","commentId":"E:AdvancedSceneManager.Core.Editor.scenesUpdated","fullName":"AdvancedSceneManager.Core.Editor.scenesUpdated","nameWithType":"Editor.scenesUpdated"},{"uid":"AdvancedSceneManager.Core.Editor.OpenSingle(UnityEditor.SceneAsset,System.Boolean)","name":"OpenSingle(SceneAsset, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_OpenSingle_UnityEditor_SceneAsset_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.OpenSingle(UnityEditor.SceneAsset,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.OpenSingle(UnityEditor.SceneAsset, System.Boolean)","nameWithType":"Editor.OpenSingle(SceneAsset, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.OpenSingle(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"OpenSingle(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_OpenSingle_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.OpenSingle(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.OpenSingle(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"Editor.OpenSingle(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"Open(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Open_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"Editor.Open(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.SceneCollection)","name":"IsOpen(SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_IsOpen_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"Editor.IsOpen(SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Editor.CanClose(AdvancedSceneManager.Models.SceneCollection)","name":"CanClose(SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_CanClose_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Editor.CanClose(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Editor.CanClose(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"Editor.CanClose(SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean,System.Boolean)","name":"Open(SceneCollection, Boolean, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Open_AdvancedSceneManager_Models_SceneCollection_System_Boolean_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.Open(AdvancedSceneManager.Models.SceneCollection, System.Boolean, System.Boolean, System.Boolean)","nameWithType":"Editor.Open(SceneCollection, Boolean, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"Close(SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Close_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"Editor.Close(SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"Close(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Close_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.Close(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"Editor.Close(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.Close(UnityEngine.SceneManagement.Scene,System.Boolean)","name":"Close(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Close_UnityEngine_SceneManagement_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.Close(UnityEngine.SceneManagement.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.Close(UnityEngine.SceneManagement.Scene, System.Boolean)","nameWithType":"Editor.Close(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.CloseAll(System.Boolean)","name":"CloseAll(Boolean)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_CloseAll_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Editor.CloseAll(System.Boolean)","fullName":"AdvancedSceneManager.Core.Editor.CloseAll(System.Boolean)","nameWithType":"Editor.CloseAll(Boolean)"},{"uid":"AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.Scene)","name":"IsOpen(Scene)","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_IsOpen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.Editor.IsOpen(AdvancedSceneManager.Models.Scene)","nameWithType":"Editor.IsOpen(Scene)"},{"uid":"AdvancedSceneManager.Core.Editor.OpenSingle*","name":"OpenSingle","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_OpenSingle_","commentId":"Overload:AdvancedSceneManager.Core.Editor.OpenSingle","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.OpenSingle","nameWithType":"Editor.OpenSingle"},{"uid":"AdvancedSceneManager.Core.Editor.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Open_","commentId":"Overload:AdvancedSceneManager.Core.Editor.Open","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.Open","nameWithType":"Editor.Open"},{"uid":"AdvancedSceneManager.Core.Editor.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_IsOpen_","commentId":"Overload:AdvancedSceneManager.Core.Editor.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.IsOpen","nameWithType":"Editor.IsOpen"},{"uid":"AdvancedSceneManager.Core.Editor.CanClose*","name":"CanClose","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_CanClose_","commentId":"Overload:AdvancedSceneManager.Core.Editor.CanClose","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.CanClose","nameWithType":"Editor.CanClose"},{"uid":"AdvancedSceneManager.Core.Editor.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_Close_","commentId":"Overload:AdvancedSceneManager.Core.Editor.Close","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.Close","nameWithType":"Editor.Close"},{"uid":"AdvancedSceneManager.Core.Editor.CloseAll*","name":"CloseAll","href":"~/api/AdvancedSceneManager.Core.Editor.yml#AdvancedSceneManager_Core_Editor_CloseAll_","commentId":"Overload:AdvancedSceneManager.Core.Editor.CloseAll","isSpec":"True","fullName":"AdvancedSceneManager.Core.Editor.CloseAll","nameWithType":"Editor.CloseAll"}],"api/AdvancedSceneManager.Core.UtilitySceneManager.yml":[{"uid":"AdvancedSceneManager.Core.UtilitySceneManager","name":"UtilitySceneManager","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml","commentId":"T:AdvancedSceneManager.Core.UtilitySceneManager","fullName":"AdvancedSceneManager.Core.UtilitySceneManager","nameWithType":"UtilitySceneManager"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.openScenes","name":"openScenes","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_openScenes","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.openScenes","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.openScenes","nameWithType":"UtilitySceneManager.openScenes"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback``1(System.Func{``0,System.Collections.IEnumerator})","name":"DoSceneCallback<T>(Func<T, IEnumerator>)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_DoSceneCallback__1_System_Func___0_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback``1(System.Func{``0,System.Collections.IEnumerator})","name.vb":"DoSceneCallback(Of T)(Func(Of T, IEnumerator))","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback<T>(System.Func<T, System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback(Of T)(System.Func(Of T, System.Collections.IEnumerator))","nameWithType":"UtilitySceneManager.DoSceneCallback<T>(Func<T, IEnumerator>)","nameWithType.vb":"UtilitySceneManager.DoSceneCallback(Of T)(Func(Of T, IEnumerator))"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.queueEmpty","name":"queueEmpty","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_queueEmpty","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.queueEmpty","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.queueEmpty","nameWithType":"UtilitySceneManager.queueEmpty"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.isBusy","name":"isBusy","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_isBusy","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.isBusy","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.isBusy","nameWithType":"UtilitySceneManager.isBusy"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.runningOperations","name":"runningOperations","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_runningOperations","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.runningOperations","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.runningOperations","nameWithType":"UtilitySceneManager.runningOperations"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations","name":"queuedOperations","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_queuedOperations","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations","nameWithType":"UtilitySceneManager.queuedOperations"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.currentOperation","name":"currentOperation","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_currentOperation","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.currentOperation","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.currentOperation","nameWithType":"UtilitySceneManager.currentOperation"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChanged","name":"ActiveSceneChanged","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_ActiveSceneChanged","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChanged","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChanged","nameWithType":"UtilitySceneManager.ActiveSceneChanged"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.SceneOpened","name":"SceneOpened","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_SceneOpened","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.SceneOpened","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.SceneOpened","nameWithType":"UtilitySceneManager.SceneOpened"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.SceneClosed","name":"SceneClosed","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_SceneClosed","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.SceneClosed","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.SceneClosed","nameWithType":"UtilitySceneManager.SceneClosed"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpening","name":"LoadingScreenOpening","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_LoadingScreenOpening","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpening","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpening","nameWithType":"UtilitySceneManager.LoadingScreenOpening"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpened","name":"LoadingScreenOpened","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_LoadingScreenOpened","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpened","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenOpened","nameWithType":"UtilitySceneManager.LoadingScreenOpened"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosing","name":"LoadingScreenClosing","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_LoadingScreenClosing","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosing","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosing","nameWithType":"UtilitySceneManager.LoadingScreenClosing"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosed","name":"LoadingScreenClosed","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_LoadingScreenClosed","commentId":"E:AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosed","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.LoadingScreenClosed","nameWithType":"UtilitySceneManager.LoadingScreenClosed"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback``1(``0,System.Action,System.Action,System.Boolean)","name":"RegisterOpenCallback<T>(T, Action, Action, Boolean)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_RegisterOpenCallback__1___0_System_Action_System_Action_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback``1(``0,System.Action,System.Action,System.Boolean)","name.vb":"RegisterOpenCallback(Of T)(T, Action, Action, Boolean)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback<T>(T, System.Action, System.Action, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback(Of T)(T, System.Action, System.Action, System.Boolean)","nameWithType":"UtilitySceneManager.RegisterOpenCallback<T>(T, Action, Action, Boolean)","nameWithType.vb":"UtilitySceneManager.RegisterOpenCallback(Of T)(T, Action, Action, Boolean)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback``1(``0,System.Action,System.Action)","name":"UnregisterCallback<T>(T, Action, Action)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_UnregisterCallback__1___0_System_Action_System_Action_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback``1(``0,System.Action,System.Action)","name.vb":"UnregisterCallback(Of T)(T, Action, Action)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback<T>(T, System.Action, System.Action)","fullName.vb":"AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback(Of T)(T, System.Action, System.Action)","nameWithType":"UtilitySceneManager.UnregisterCallback<T>(T, Action, Action)","nameWithType.vb":"UtilitySceneManager.UnregisterCallback(Of T)(T, Action, Action)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Reopen(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Reopen(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Reopen_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.Reopen(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Reopen(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"UtilitySceneManager.Reopen(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","name":"OpenOrReopen(Scene, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_OpenOrReopen_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"UtilitySceneManager.OpenOrReopen(Scene, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Close(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Close_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Close(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"UtilitySceneManager.Close(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.CloseAll(System.Boolean)","name":"CloseAll(Boolean)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_CloseAll_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.CloseAll(System.Boolean)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.CloseAll(System.Boolean)","nameWithType":"UtilitySceneManager.CloseAll(Boolean)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(AdvancedSceneManager.Models.Scene,System.Nullable{System.Boolean})","name":"Toggle(Scene, Nullable<Boolean>)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Toggle_AdvancedSceneManager_Models_Scene_System_Nullable_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.Toggle(AdvancedSceneManager.Models.Scene,System.Nullable{System.Boolean})","name.vb":"Toggle(Scene, Nullable(Of Boolean))","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(AdvancedSceneManager.Models.Scene, System.Nullable<System.Boolean>)","fullName.vb":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(AdvancedSceneManager.Models.Scene, System.Nullable(Of System.Boolean))","nameWithType":"UtilitySceneManager.Toggle(Scene, Nullable<Boolean>)","nameWithType.vb":"UtilitySceneManager.Toggle(Scene, Nullable(Of Boolean))"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(UnityEngine.SceneManagement.Scene,System.Nullable{System.Boolean})","name":"Toggle(Scene, Nullable<Boolean>)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Toggle_UnityEngine_SceneManagement_Scene_System_Nullable_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.Toggle(UnityEngine.SceneManagement.Scene,System.Nullable{System.Boolean})","name.vb":"Toggle(Scene, Nullable(Of Boolean))","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(UnityEngine.SceneManagement.Scene, System.Nullable<System.Boolean>)","fullName.vb":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle(UnityEngine.SceneManagement.Scene, System.Nullable(Of System.Boolean))","nameWithType":"UtilitySceneManager.Toggle(Scene, Nullable<Boolean>)","nameWithType.vb":"UtilitySceneManager.Toggle(Scene, Nullable(Of Boolean))"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(AdvancedSceneManager.Models.Scene)","name":"IsOpen(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_IsOpen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(AdvancedSceneManager.Models.Scene)","nameWithType":"UtilitySceneManager.IsOpen(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(UnityEngine.SceneManagement.Scene)","name":"IsOpen(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_IsOpen_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen(UnityEngine.SceneManagement.Scene)","nameWithType":"UtilitySceneManager.IsOpen(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(UnityEngine.SceneManagement.Scene)","name":"FindOpenScene(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindOpenScene_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(UnityEngine.SceneManagement.Scene)","nameWithType":"UtilitySceneManager.FindOpenScene(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(AdvancedSceneManager.Models.Scene)","name":"FindOpenScene(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindOpenScene_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene(AdvancedSceneManager.Models.Scene)","nameWithType":"UtilitySceneManager.FindOpenScene(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(AdvancedSceneManager.Models.Scene)","name":"FindPreloadedScene(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindPreloadedScene_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(AdvancedSceneManager.Models.Scene)","nameWithType":"UtilitySceneManager.FindPreloadedScene(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(UnityEngine.SceneManagement.Scene)","name":"FindPreloadedScene(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindPreloadedScene_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene(UnityEngine.SceneManagement.Scene)","nameWithType":"UtilitySceneManager.FindPreloadedScene(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes","name":"FindPreloadedScenes()","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindPreloadedScenes","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes()","nameWithType":"UtilitySceneManager.FindPreloadedScenes()"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive(UnityEngine.SceneManagement.Scene)","name":"SetActive(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_SetActive_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.SetActive(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive(UnityEngine.SceneManagement.Scene)","nameWithType":"UtilitySceneManager.SetActive(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive(AdvancedSceneManager.Models.Scene)","name":"SetActive(Scene)","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_SetActive_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.UtilitySceneManager.SetActive(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive(AdvancedSceneManager.Models.Scene)","nameWithType":"UtilitySceneManager.SetActive(Scene)"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.activeScene","name":"activeScene","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_activeScene","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.activeScene","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.activeScene","nameWithType":"UtilitySceneManager.activeScene"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad","name":"dontDestroyOnLoad","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_dontDestroyOnLoad","commentId":"P:AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad","nameWithType":"UtilitySceneManager.dontDestroyOnLoad"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.openScenes*","name":"openScenes","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_openScenes_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.openScenes","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.openScenes","nameWithType":"UtilitySceneManager.openScenes"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback*","name":"DoSceneCallback","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_DoSceneCallback_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.DoSceneCallback","nameWithType":"UtilitySceneManager.DoSceneCallback"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.isBusy*","name":"isBusy","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_isBusy_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.isBusy","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.isBusy","nameWithType":"UtilitySceneManager.isBusy"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.runningOperations*","name":"runningOperations","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_runningOperations_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.runningOperations","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.runningOperations","nameWithType":"UtilitySceneManager.runningOperations"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations*","name":"queuedOperations","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_queuedOperations_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.queuedOperations","nameWithType":"UtilitySceneManager.queuedOperations"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.currentOperation*","name":"currentOperation","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_currentOperation_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.currentOperation","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.currentOperation","nameWithType":"UtilitySceneManager.currentOperation"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback*","name":"RegisterOpenCallback","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_RegisterOpenCallback_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.RegisterOpenCallback","nameWithType":"UtilitySceneManager.RegisterOpenCallback"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback*","name":"UnregisterCallback","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_UnregisterCallback_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.UnregisterCallback","nameWithType":"UtilitySceneManager.UnregisterCallback"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Reopen_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Reopen","nameWithType":"UtilitySceneManager.Reopen"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen*","name":"OpenOrReopen","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_OpenOrReopen_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.OpenOrReopen","nameWithType":"UtilitySceneManager.OpenOrReopen"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Close_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.Close","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Close","nameWithType":"UtilitySceneManager.Close"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.CloseAll*","name":"CloseAll","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_CloseAll_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.CloseAll","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.CloseAll","nameWithType":"UtilitySceneManager.CloseAll"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_Toggle_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.Toggle","nameWithType":"UtilitySceneManager.Toggle"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_IsOpen_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.IsOpen","nameWithType":"UtilitySceneManager.IsOpen"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene*","name":"FindOpenScene","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindOpenScene_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindOpenScene","nameWithType":"UtilitySceneManager.FindOpenScene"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene*","name":"FindPreloadedScene","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindPreloadedScene_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScene","nameWithType":"UtilitySceneManager.FindPreloadedScene"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes*","name":"FindPreloadedScenes","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_FindPreloadedScenes_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.FindPreloadedScenes","nameWithType":"UtilitySceneManager.FindPreloadedScenes"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive*","name":"SetActive","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_SetActive_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.SetActive","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.SetActive","nameWithType":"UtilitySceneManager.SetActive"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.activeScene*","name":"activeScene","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_activeScene_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.activeScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.activeScene","nameWithType":"UtilitySceneManager.activeScene"},{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad*","name":"dontDestroyOnLoad","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.yml#AdvancedSceneManager_Core_UtilitySceneManager_dontDestroyOnLoad_","commentId":"Overload:AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad","isSpec":"True","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.dontDestroyOnLoad","nameWithType":"UtilitySceneManager.dontDestroyOnLoad"}],"api/AdvancedSceneManager.Core.yml":[{"uid":"AdvancedSceneManager.Core","name":"AdvancedSceneManager.Core","href":"~/api/AdvancedSceneManager.Core.yml","commentId":"N:AdvancedSceneManager.Core","fullName":"AdvancedSceneManager.Core","nameWithType":"AdvancedSceneManager.Core"}],"api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml":[{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1","name":"EditorWindow_UIElements<T>","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml","commentId":"T:AdvancedSceneManager.Editor.EditorWindow_UIElements`1","name.vb":"EditorWindow_UIElements(Of T)","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T)","nameWithType":"EditorWindow_UIElements<T>","nameWithType.vb":"EditorWindow_UIElements(Of T)"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.autoReloadOnWindowFocus","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_autoReloadOnWindowFocus","commentId":"P:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.autoReloadOnWindowFocus","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.autoReloadOnWindowFocus","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).autoReloadOnWindowFocus","nameWithType":"EditorWindow_UIElements<T>.autoReloadOnWindowFocus","nameWithType.vb":"EditorWindow_UIElements(Of T).autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_path","commentId":"P:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.path","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.path","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).path","nameWithType":"EditorWindow_UIElements<T>.path","nameWithType.vb":"EditorWindow_UIElements(Of T).path"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_title","commentId":"P:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.title","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.title","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).title","nameWithType":"EditorWindow_UIElements<T>.title","nameWithType.vb":"EditorWindow_UIElements(Of T).title"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.window","name":"window","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_window","commentId":"P:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.window","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.window","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).window","nameWithType":"EditorWindow_UIElements<T>.window","nameWithType.vb":"EditorWindow_UIElements(Of T).window"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Open","name":"Open()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Open","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Open","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Open()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Open()","nameWithType":"EditorWindow_UIElements<T>.Open()","nameWithType.vb":"EditorWindow_UIElements(Of T).Open()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Close","name":"Close()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Close","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Close","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Close()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Close()","nameWithType":"EditorWindow_UIElements<T>.Close()","nameWithType.vb":"EditorWindow_UIElements(Of T).Close()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnClose","name":"OnClose()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnClose","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnClose","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnClose()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnClose()","nameWithType":"EditorWindow_UIElements<T>.OnClose()","nameWithType.vb":"EditorWindow_UIElements(Of T).OnClose()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.DoShow","name":"DoShow()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_DoShow","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.DoShow","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.DoShow()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).DoShow()","nameWithType":"EditorWindow_UIElements<T>.DoShow()","nameWithType.vb":"EditorWindow_UIElements(Of T).DoShow()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnShow","name":"OnShow()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnShow","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnShow","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnShow()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnShow()","nameWithType":"EditorWindow_UIElements<T>.OnShow()","nameWithType.vb":"EditorWindow_UIElements(Of T).OnShow()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Reopen","name":"Reopen()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Reopen","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Reopen","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Reopen()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Reopen()","nameWithType":"EditorWindow_UIElements<T>.Reopen()","nameWithType.vb":"EditorWindow_UIElements(Of T).Reopen()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.isMainContentLoaded","name":"isMainContentLoaded","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_isMainContentLoaded","commentId":"P:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.isMainContentLoaded","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.isMainContentLoaded","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).isMainContentLoaded","nameWithType":"EditorWindow_UIElements<T>.isMainContentLoaded","nameWithType.vb":"EditorWindow_UIElements(Of T).isMainContentLoaded"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ShowSuspendMessage","name":"ShowSuspendMessage()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_ShowSuspendMessage","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ShowSuspendMessage","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.ShowSuspendMessage()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).ShowSuspendMessage()","nameWithType":"EditorWindow_UIElements<T>.ShowSuspendMessage()","nameWithType.vb":"EditorWindow_UIElements(Of T).ShowSuspendMessage()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement)","name":"LoadContent(String, VisualElement)","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_LoadContent_System_String_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.LoadContent(System.String, UnityEngine.UIElements.VisualElement)","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).LoadContent(System.String, UnityEngine.UIElements.VisualElement)","nameWithType":"EditorWindow_UIElements<T>.LoadContent(String, VisualElement)","nameWithType.vb":"EditorWindow_UIElements(Of T).LoadContent(String, VisualElement)"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement,System.Boolean,System.Boolean,System.Boolean)","name":"LoadContent(String, VisualElement, Boolean, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_LoadContent_System_String_UnityEngine_UIElements_VisualElement_System_Boolean_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement,System.Boolean,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.LoadContent(System.String, UnityEngine.UIElements.VisualElement, System.Boolean, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).LoadContent(System.String, UnityEngine.UIElements.VisualElement, System.Boolean, System.Boolean, System.Boolean)","nameWithType":"EditorWindow_UIElements<T>.LoadContent(String, VisualElement, Boolean, Boolean, Boolean)","nameWithType.vb":"EditorWindow_UIElements(Of T).LoadContent(String, VisualElement, Boolean, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ReloadContent","name":"ReloadContent()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_ReloadContent","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ReloadContent","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.ReloadContent()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).ReloadContent()","nameWithType":"EditorWindow_UIElements<T>.ReloadContent()","nameWithType.vb":"EditorWindow_UIElements(Of T).ReloadContent()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnFocus","name":"OnFocus()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnFocus","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnFocus","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnFocus()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnFocus()","nameWithType":"EditorWindow_UIElements<T>.OnFocus()","nameWithType.vb":"EditorWindow_UIElements(Of T).OnFocus()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnEnable","name":"OnEnable()","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnEnable","commentId":"M:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnEnable","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnEnable()","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnEnable()","nameWithType":"EditorWindow_UIElements<T>.OnEnable()","nameWithType.vb":"EditorWindow_UIElements(Of T).OnEnable()"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.autoReloadOnWindowFocus*","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_autoReloadOnWindowFocus_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.autoReloadOnWindowFocus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.autoReloadOnWindowFocus","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).autoReloadOnWindowFocus","nameWithType":"EditorWindow_UIElements<T>.autoReloadOnWindowFocus","nameWithType.vb":"EditorWindow_UIElements(Of T).autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_path_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.path","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).path","nameWithType":"EditorWindow_UIElements<T>.path","nameWithType.vb":"EditorWindow_UIElements(Of T).path"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_title_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.title","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).title","nameWithType":"EditorWindow_UIElements<T>.title","nameWithType.vb":"EditorWindow_UIElements(Of T).title"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.window*","name":"window","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_window_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.window","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.window","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).window","nameWithType":"EditorWindow_UIElements<T>.window","nameWithType.vb":"EditorWindow_UIElements(Of T).window"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Open_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Open","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Open","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Open","nameWithType":"EditorWindow_UIElements<T>.Open","nameWithType.vb":"EditorWindow_UIElements(Of T).Open"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Close_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Close","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Close","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Close","nameWithType":"EditorWindow_UIElements<T>.Close","nameWithType.vb":"EditorWindow_UIElements(Of T).Close"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnClose_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnClose","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnClose","nameWithType":"EditorWindow_UIElements<T>.OnClose","nameWithType.vb":"EditorWindow_UIElements(Of T).OnClose"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.DoShow*","name":"DoShow","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_DoShow_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.DoShow","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.DoShow","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).DoShow","nameWithType":"EditorWindow_UIElements<T>.DoShow","nameWithType.vb":"EditorWindow_UIElements(Of T).DoShow"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnShow*","name":"OnShow","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnShow_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnShow","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnShow","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnShow","nameWithType":"EditorWindow_UIElements<T>.OnShow","nameWithType.vb":"EditorWindow_UIElements(Of T).OnShow"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_Reopen_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.Reopen","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).Reopen","nameWithType":"EditorWindow_UIElements<T>.Reopen","nameWithType.vb":"EditorWindow_UIElements(Of T).Reopen"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.isMainContentLoaded*","name":"isMainContentLoaded","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_isMainContentLoaded_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.isMainContentLoaded","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.isMainContentLoaded","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).isMainContentLoaded","nameWithType":"EditorWindow_UIElements<T>.isMainContentLoaded","nameWithType.vb":"EditorWindow_UIElements(Of T).isMainContentLoaded"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ShowSuspendMessage*","name":"ShowSuspendMessage","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_ShowSuspendMessage_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ShowSuspendMessage","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.ShowSuspendMessage","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).ShowSuspendMessage","nameWithType":"EditorWindow_UIElements<T>.ShowSuspendMessage","nameWithType.vb":"EditorWindow_UIElements(Of T).ShowSuspendMessage"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent*","name":"LoadContent","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_LoadContent_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.LoadContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.LoadContent","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).LoadContent","nameWithType":"EditorWindow_UIElements<T>.LoadContent","nameWithType.vb":"EditorWindow_UIElements(Of T).LoadContent"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ReloadContent*","name":"ReloadContent","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_ReloadContent_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.ReloadContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.ReloadContent","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).ReloadContent","nameWithType":"EditorWindow_UIElements<T>.ReloadContent","nameWithType.vb":"EditorWindow_UIElements(Of T).ReloadContent"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnFocus*","name":"OnFocus","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnFocus_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnFocus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnFocus","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnFocus","nameWithType":"EditorWindow_UIElements<T>.OnFocus","nameWithType.vb":"EditorWindow_UIElements(Of T).OnFocus"},{"uid":"AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.EditorWindow_UIElements-1.yml#AdvancedSceneManager_Editor_EditorWindow_UIElements_1_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.EditorWindow_UIElements`1.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditorWindow_UIElements<T>.OnEnable","fullName.vb":"AdvancedSceneManager.Editor.EditorWindow_UIElements(Of T).OnEnable","nameWithType":"EditorWindow_UIElements<T>.OnEnable","nameWithType.vb":"EditorWindow_UIElements(Of T).OnEnable"}],"api/AdvancedSceneManager.Editor.GenericPopup.Item.yml":[{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item","name":"GenericPopup.Item","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml","commentId":"T:AdvancedSceneManager.Editor.GenericPopup.Item","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item","nameWithType":"GenericPopup.Item"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.Separator","name":"Separator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_Separator","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.Separator","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.Separator","nameWithType":"GenericPopup.Item.Separator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.name","name":"name","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_name","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.name","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.name","nameWithType":"GenericPopup.Item.name"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isChecked","name":"isChecked","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isChecked","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isChecked","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isChecked","nameWithType":"GenericPopup.Item.isChecked"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.onClick","name":"onClick","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_onClick","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.onClick","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.onClick","nameWithType":"GenericPopup.Item.onClick"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable","name":"isCheckable","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isCheckable","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable","nameWithType":"GenericPopup.Item.isCheckable"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled","name":"isEnabled","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isEnabled","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled","nameWithType":"GenericPopup.Item.isEnabled"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isVisible","name":"isVisible","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isVisible","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isVisible","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isVisible","nameWithType":"GenericPopup.Item.isVisible"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isBold","name":"isBold","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isBold","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isBold","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isBold","nameWithType":"GenericPopup.Item.isBold"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator","name":"isSeparator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isSeparator","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator","nameWithType":"GenericPopup.Item.isSeparator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String)","name":"Create(String)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_Create_System_String_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String)","nameWithType":"GenericPopup.Item.Create(String)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String,System.Action)","name":"Create(String, Action)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_Create_System_String_System_Action_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String,System.Action)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.Create(System.String, System.Action)","nameWithType":"GenericPopup.Item.Create(String, Action)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable","name":"AsCheckable()","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_AsCheckable","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable()","nameWithType":"GenericPopup.Item.AsCheckable()"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable(System.Action{System.Boolean})","name":"AsCheckable(Action<Boolean>)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_AsCheckable_System_Action_System_Boolean__","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable(System.Action{System.Boolean})","name.vb":"AsCheckable(Action(Of Boolean))","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable(System.Action<System.Boolean>)","fullName.vb":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable(System.Action(Of System.Boolean))","nameWithType":"GenericPopup.Item.AsCheckable(Action<Boolean>)","nameWithType.vb":"GenericPopup.Item.AsCheckable(Action(Of Boolean))"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus(System.Boolean)","name":"WithCheckedStatus(Boolean)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithCheckedStatus_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus(System.Boolean)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus(System.Boolean)","nameWithType":"GenericPopup.Item.WithCheckedStatus(Boolean)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState(System.Boolean)","name":"WithEnabledState(Boolean)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithEnabledState_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState(System.Boolean)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState(System.Boolean)","nameWithType":"GenericPopup.Item.WithEnabledState(Boolean)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked(System.Action)","name":"WhenClicked(Action)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WhenClicked_System_Action_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked(System.Action)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked(System.Action)","nameWithType":"GenericPopup.Item.WhenClicked(Action)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState(System.Boolean)","name":"WithVisibleState(Boolean)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithVisibleState_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState(System.Boolean)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState(System.Boolean)","nameWithType":"GenericPopup.Item.WithVisibleState(Boolean)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState(System.Boolean)","name":"WithBoldState(Boolean)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithBoldState_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState(System.Boolean)","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState(System.Boolean)","nameWithType":"GenericPopup.Item.WithBoldState(Boolean)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.Separator*","name":"Separator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_Separator_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.Separator","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.Separator","nameWithType":"GenericPopup.Item.Separator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.name*","name":"name","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_name_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.name","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.name","nameWithType":"GenericPopup.Item.name"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isChecked*","name":"isChecked","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isChecked_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isChecked","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isChecked","nameWithType":"GenericPopup.Item.isChecked"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.onClick*","name":"onClick","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_onClick_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.onClick","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.onClick","nameWithType":"GenericPopup.Item.onClick"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable*","name":"isCheckable","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isCheckable_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isCheckable","nameWithType":"GenericPopup.Item.isCheckable"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled*","name":"isEnabled","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isEnabled_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isEnabled","nameWithType":"GenericPopup.Item.isEnabled"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isVisible*","name":"isVisible","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isVisible_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isVisible","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isVisible","nameWithType":"GenericPopup.Item.isVisible"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isBold*","name":"isBold","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isBold_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isBold","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isBold","nameWithType":"GenericPopup.Item.isBold"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator*","name":"isSeparator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_isSeparator_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.isSeparator","nameWithType":"GenericPopup.Item.isSeparator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.Create*","name":"Create","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_Create_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.Create","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.Create","nameWithType":"GenericPopup.Item.Create"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable*","name":"AsCheckable","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_AsCheckable_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.AsCheckable","nameWithType":"GenericPopup.Item.AsCheckable"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus*","name":"WithCheckedStatus","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithCheckedStatus_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithCheckedStatus","nameWithType":"GenericPopup.Item.WithCheckedStatus"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState*","name":"WithEnabledState","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithEnabledState_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithEnabledState","nameWithType":"GenericPopup.Item.WithEnabledState"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked*","name":"WhenClicked","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WhenClicked_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WhenClicked","nameWithType":"GenericPopup.Item.WhenClicked"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState*","name":"WithVisibleState","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithVisibleState_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithVisibleState","nameWithType":"GenericPopup.Item.WithVisibleState"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState*","name":"WithBoldState","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.Item.yml#AdvancedSceneManager_Editor_GenericPopup_Item_WithBoldState_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Item.WithBoldState","nameWithType":"GenericPopup.Item.WithBoldState"}],"api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml":[{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup","name":"OpenInEditorPopup","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml","commentId":"T:AdvancedSceneManager.Editor.OpenInEditorPopup","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup","nameWithType":"OpenInEditorPopup"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_path","commentId":"P:AdvancedSceneManager.Editor.OpenInEditorPopup.path","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.path","nameWithType":"OpenInEditorPopup.path"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.height","name":"height","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_height","commentId":"P:AdvancedSceneManager.Editor.OpenInEditorPopup.height","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.height","nameWithType":"OpenInEditorPopup.height"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh(AdvancedSceneManager.Models.Scene)","name":"Refresh(Scene)","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_Refresh_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh(AdvancedSceneManager.Models.Scene)","nameWithType":"OpenInEditorPopup.Refresh(Scene)"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen(AdvancedSceneManager.Editor.OpenInEditorPopup)","name":"OnReopen(OpenInEditorPopup)","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_OnReopen_AdvancedSceneManager_Editor_OpenInEditorPopup_","commentId":"M:AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen(AdvancedSceneManager.Editor.OpenInEditorPopup)","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen(AdvancedSceneManager.Editor.OpenInEditorPopup)","nameWithType":"OpenInEditorPopup.OnReopen(OpenInEditorPopup)"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_path_","commentId":"Overload:AdvancedSceneManager.Editor.OpenInEditorPopup.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.path","nameWithType":"OpenInEditorPopup.path"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.height*","name":"height","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_height_","commentId":"Overload:AdvancedSceneManager.Editor.OpenInEditorPopup.height","isSpec":"True","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.height","nameWithType":"OpenInEditorPopup.height"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh*","name":"Refresh","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_Refresh_","commentId":"Overload:AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.Refresh","nameWithType":"OpenInEditorPopup.Refresh"},{"uid":"AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen*","name":"OnReopen","href":"~/api/AdvancedSceneManager.Editor.OpenInEditorPopup.yml#AdvancedSceneManager_Editor_OpenInEditorPopup_OnReopen_","commentId":"Overload:AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.OpenInEditorPopup.OnReopen","nameWithType":"OpenInEditorPopup.OnReopen"}],"api/AdvancedSceneManager.Editor.PickTagPopup.yml":[{"uid":"AdvancedSceneManager.Editor.PickTagPopup","name":"PickTagPopup","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml","commentId":"T:AdvancedSceneManager.Editor.PickTagPopup","fullName":"AdvancedSceneManager.Editor.PickTagPopup","nameWithType":"PickTagPopup"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_path","commentId":"P:AdvancedSceneManager.Editor.PickTagPopup.path","fullName":"AdvancedSceneManager.Editor.PickTagPopup.path","nameWithType":"PickTagPopup.path"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.enableBorder","name":"enableBorder","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_enableBorder","commentId":"P:AdvancedSceneManager.Editor.PickTagPopup.enableBorder","fullName":"AdvancedSceneManager.Editor.PickTagPopup.enableBorder","nameWithType":"PickTagPopup.enableBorder"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.Refresh(AdvancedSceneManager.Models.SceneTag,System.Action{AdvancedSceneManager.Models.SceneTag})","name":"Refresh(SceneTag, Action<SceneTag>)","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_Refresh_AdvancedSceneManager_Models_SceneTag_System_Action_AdvancedSceneManager_Models_SceneTag__","commentId":"M:AdvancedSceneManager.Editor.PickTagPopup.Refresh(AdvancedSceneManager.Models.SceneTag,System.Action{AdvancedSceneManager.Models.SceneTag})","name.vb":"Refresh(SceneTag, Action(Of SceneTag))","fullName":"AdvancedSceneManager.Editor.PickTagPopup.Refresh(AdvancedSceneManager.Models.SceneTag, System.Action<AdvancedSceneManager.Models.SceneTag>)","fullName.vb":"AdvancedSceneManager.Editor.PickTagPopup.Refresh(AdvancedSceneManager.Models.SceneTag, System.Action(Of AdvancedSceneManager.Models.SceneTag))","nameWithType":"PickTagPopup.Refresh(SceneTag, Action<SceneTag>)","nameWithType.vb":"PickTagPopup.Refresh(SceneTag, Action(Of SceneTag))"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.OnReopen(AdvancedSceneManager.Editor.PickTagPopup)","name":"OnReopen(PickTagPopup)","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_OnReopen_AdvancedSceneManager_Editor_PickTagPopup_","commentId":"M:AdvancedSceneManager.Editor.PickTagPopup.OnReopen(AdvancedSceneManager.Editor.PickTagPopup)","fullName":"AdvancedSceneManager.Editor.PickTagPopup.OnReopen(AdvancedSceneManager.Editor.PickTagPopup)","nameWithType":"PickTagPopup.OnReopen(PickTagPopup)"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_path_","commentId":"Overload:AdvancedSceneManager.Editor.PickTagPopup.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.PickTagPopup.path","nameWithType":"PickTagPopup.path"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.enableBorder*","name":"enableBorder","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_enableBorder_","commentId":"Overload:AdvancedSceneManager.Editor.PickTagPopup.enableBorder","isSpec":"True","fullName":"AdvancedSceneManager.Editor.PickTagPopup.enableBorder","nameWithType":"PickTagPopup.enableBorder"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.Refresh*","name":"Refresh","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_Refresh_","commentId":"Overload:AdvancedSceneManager.Editor.PickTagPopup.Refresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.PickTagPopup.Refresh","nameWithType":"PickTagPopup.Refresh"},{"uid":"AdvancedSceneManager.Editor.PickTagPopup.OnReopen*","name":"OnReopen","href":"~/api/AdvancedSceneManager.Editor.PickTagPopup.yml#AdvancedSceneManager_Editor_PickTagPopup_OnReopen_","commentId":"Overload:AdvancedSceneManager.Editor.PickTagPopup.OnReopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.PickTagPopup.OnReopen","nameWithType":"PickTagPopup.OnReopen"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.Tab.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab","name":"SceneManagerWindow.Tab","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.Tab.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow.Tab","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab","nameWithType":"SceneManagerWindow.Tab"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Scenes","name":"Scenes","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.Tab.yml#AdvancedSceneManager_Editor_SceneManagerWindow_Tab_Scenes","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Scenes","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Scenes","nameWithType":"SceneManagerWindow.Tab.Scenes"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Tags","name":"Tags","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.Tab.yml#AdvancedSceneManager_Editor_SceneManagerWindow_Tab_Tags","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Tags","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Tags","nameWithType":"SceneManagerWindow.Tab.Tags"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Settings","name":"Settings","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.Tab.yml#AdvancedSceneManager_Editor_SceneManagerWindow_Tab_Settings","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Settings","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Tab.Settings","nameWithType":"SceneManagerWindow.Tab.Settings"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow","name":"SceneManagerWindow","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow","nameWithType":"SceneManagerWindow"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.OnGUIEvent","name":"OnGUIEvent","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_OnGUIEvent","commentId":"E:AdvancedSceneManager.Editor.SceneManagerWindow.OnGUIEvent","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.OnGUIEvent","nameWithType":"SceneManagerWindow.OnGUIEvent"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.MouseUp","name":"MouseUp","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_MouseUp","commentId":"E:AdvancedSceneManager.Editor.SceneManagerWindow.MouseUp","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.MouseUp","nameWithType":"SceneManagerWindow.MouseUp"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.position","name":"position","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_position","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.position","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.position","nameWithType":"SceneManagerWindow.position"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode","name":"IsDarkMode","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_IsDarkMode","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode","nameWithType":"SceneManagerWindow.IsDarkMode"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_path","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.path","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.path","nameWithType":"SceneManagerWindow.path"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_autoReloadOnWindowFocus","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus","nameWithType":"SceneManagerWindow.autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged","name":"IgnoreProfileChanged()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_IgnoreProfileChanged","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged()","nameWithType":"SceneManagerWindow.IgnoreProfileChanged()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable","name":"OnEnable()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_OnEnable","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable()","nameWithType":"SceneManagerWindow.OnEnable()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage","name":"deleteTempBuildMessage","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_deleteTempBuildMessage","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage","nameWithType":"SceneManagerWindow.deleteTempBuildMessage"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus","name":"OnFocus()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_OnFocus","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus()","nameWithType":"SceneManagerWindow.OnFocus()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab","name":"ReopenTab()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_ReopenTab","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab()","nameWithType":"SceneManagerWindow.ReopenTab()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Save(UnityEngine.ScriptableObject,System.Boolean)","name":"Save(ScriptableObject, Boolean)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_Save_UnityEngine_ScriptableObject_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.Save(UnityEngine.ScriptableObject,System.Boolean)","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Save(UnityEngine.ScriptableObject, System.Boolean)","nameWithType":"SceneManagerWindow.Save(ScriptableObject, Boolean)"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode*","name":"IsDarkMode","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_IsDarkMode_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.IsDarkMode","nameWithType":"SceneManagerWindow.IsDarkMode"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_path_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.path","nameWithType":"SceneManagerWindow.path"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus*","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_autoReloadOnWindowFocus_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.autoReloadOnWindowFocus","nameWithType":"SceneManagerWindow.autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged*","name":"IgnoreProfileChanged","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_IgnoreProfileChanged_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.IgnoreProfileChanged","nameWithType":"SceneManagerWindow.IgnoreProfileChanged"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.OnEnable","nameWithType":"SceneManagerWindow.OnEnable"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage*","name":"deleteTempBuildMessage","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_deleteTempBuildMessage_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.deleteTempBuildMessage","nameWithType":"SceneManagerWindow.deleteTempBuildMessage"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus*","name":"OnFocus","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_OnFocus_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.OnFocus","nameWithType":"SceneManagerWindow.OnFocus"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab*","name":"ReopenTab","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_ReopenTab_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.ReopenTab","nameWithType":"SceneManagerWindow.ReopenTab"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.Save*","name":"Save","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.yml#AdvancedSceneManager_Editor_SceneManagerWindow_Save_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.Save","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.Save","nameWithType":"SceneManagerWindow.Save"}],"api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility","name":"BuildSettingsUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility","nameWithType":"BuildSettingsUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings","name":"UpdateBuildSettings()","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_UpdateBuildSettings","commentId":"M:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings()","nameWithType":"BuildSettingsUtility.UpdateBuildSettings()"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList","name":"GetOrderedList()","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_GetOrderedList","commentId":"M:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList()","nameWithType":"BuildSettingsUtility.GetOrderedList()"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded(AdvancedSceneManager.Models.Scene)","name":"IsIncluded(Scene)","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_IsIncluded_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded(AdvancedSceneManager.Models.Scene)","nameWithType":"BuildSettingsUtility.IsIncluded(Scene)"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState(System.String)","name":"GetEnabledState(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_GetEnabledState_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState(System.String)","nameWithType":"BuildSettingsUtility.GetEnabledState(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings*","name":"UpdateBuildSettings","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_UpdateBuildSettings_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.UpdateBuildSettings","nameWithType":"BuildSettingsUtility.UpdateBuildSettings"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList*","name":"GetOrderedList","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_GetOrderedList_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetOrderedList","nameWithType":"BuildSettingsUtility.GetOrderedList"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded*","name":"IsIncluded","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_IsIncluded_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.IsIncluded","nameWithType":"BuildSettingsUtility.IsIncluded"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState*","name":"GetEnabledState","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_GetEnabledState_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.GetEnabledState","nameWithType":"BuildSettingsUtility.GetEnabledState"}],"api/AdvancedSceneManager.Editor.Utility.EditorFolderUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility","name":"EditorFolderUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorFolderUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.EditorFolderUtility","fullName":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility","nameWithType":"EditorFolderUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists(System.String)","name":"EnsureFolderExists(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorFolderUtility.yml#AdvancedSceneManager_Editor_Utility_EditorFolderUtility_EnsureFolderExists_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists(System.String)","nameWithType":"EditorFolderUtility.EnsureFolderExists(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists*","name":"EnsureFolderExists","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorFolderUtility.yml#AdvancedSceneManager_Editor_Utility_EditorFolderUtility_EnsureFolderExists_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.EditorFolderUtility.EnsureFolderExists","nameWithType":"EditorFolderUtility.EnsureFolderExists"}],"api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions","name":"VisualElementExtensions","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.VisualElementExtensions","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions","nameWithType":"VisualElementExtensions"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor","name":"DefaultBackgroundColor","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_DefaultBackgroundColor","commentId":"P:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor","nameWithType":"VisualElementExtensions.DefaultBackgroundColor"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt``1(``0,System.Boolean)","name":"SetEnabledExt<TElement>(TElement, Boolean)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_SetEnabledExt__1___0_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt``1(``0,System.Boolean)","name.vb":"SetEnabledExt(Of TElement)(TElement, Boolean)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt<TElement>(TElement, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt(Of TElement)(TElement, System.Boolean)","nameWithType":"VisualElementExtensions.SetEnabledExt<TElement>(TElement, Boolean)","nameWithType.vb":"VisualElementExtensions.SetEnabledExt(Of TElement)(TElement, Boolean)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt(UnityEditor.UIElements.EnumField,System.Enum)","name":"SetValueWithoutNotifyExt(EnumField, Enum)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_SetValueWithoutNotifyExt_UnityEditor_UIElements_EnumField_System_Enum_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt(UnityEditor.UIElements.EnumField,System.Enum)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt(UnityEditor.UIElements.EnumField, System.Enum)","nameWithType":"VisualElementExtensions.SetValueWithoutNotifyExt(EnumField, Enum)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup``1(AdvancedSceneManager.Editor.SceneField,System.String,``0,System.String,System.Action,System.Boolean,System.String)","name":"Setup<T>(SceneField, String, T, String, Action, Boolean, String)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_Setup__1_AdvancedSceneManager_Editor_SceneField_System_String___0_System_String_System_Action_System_Boolean_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup``1(AdvancedSceneManager.Editor.SceneField,System.String,``0,System.String,System.Action,System.Boolean,System.String)","name.vb":"Setup(Of T)(SceneField, String, T, String, Action, Boolean, String)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup<T>(AdvancedSceneManager.Editor.SceneField, System.String, T, System.String, System.Action, System.Boolean, System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(Of T)(AdvancedSceneManager.Editor.SceneField, System.String, T, System.String, System.Action, System.Boolean, System.String)","nameWithType":"VisualElementExtensions.Setup<T>(SceneField, String, T, String, Action, Boolean, String)","nameWithType.vb":"VisualElementExtensions.Setup(Of T)(SceneField, String, T, String, Action, Boolean, String)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup``2(``0,``1,System.String,System.Action,System.Boolean,System.String)","name":"Setup<TElement, T>(TElement, T, String, Action, Boolean, String)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_Setup__2___0___1_System_String_System_Action_System_Boolean_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup``2(``0,``1,System.String,System.Action,System.Boolean,System.String)","name.vb":"Setup(Of TElement, T)(TElement, T, String, Action, Boolean, String)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup<TElement, T>(TElement, T, System.String, System.Action, System.Boolean, System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(Of TElement, T)(TElement, T, System.String, System.Action, System.Boolean, System.String)","nameWithType":"VisualElementExtensions.Setup<TElement, T>(TElement, T, String, Action, Boolean, String)","nameWithType.vb":"VisualElementExtensions.Setup(Of TElement, T)(TElement, T, String, Action, Boolean, String)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Toggle,UnityEngine.UIElements.EventCallback{UnityEngine.UIElements.ChangeEvent{System.Boolean}},System.Boolean,System.String)","name":"Setup(Toggle, EventCallback<ChangeEvent<Boolean>>, Boolean, String)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_Setup_UnityEngine_UIElements_Toggle_UnityEngine_UIElements_EventCallback_UnityEngine_UIElements_ChangeEvent_System_Boolean___System_Boolean_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Toggle,UnityEngine.UIElements.EventCallback{UnityEngine.UIElements.ChangeEvent{System.Boolean}},System.Boolean,System.String)","name.vb":"Setup(Toggle, EventCallback(Of ChangeEvent(Of Boolean)), Boolean, String)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Toggle, UnityEngine.UIElements.EventCallback<UnityEngine.UIElements.ChangeEvent<System.Boolean>>, System.Boolean, System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Toggle, UnityEngine.UIElements.EventCallback(Of UnityEngine.UIElements.ChangeEvent(Of System.Boolean)), System.Boolean, System.String)","nameWithType":"VisualElementExtensions.Setup(Toggle, EventCallback<ChangeEvent<Boolean>>, Boolean, String)","nameWithType.vb":"VisualElementExtensions.Setup(Toggle, EventCallback(Of ChangeEvent(Of Boolean)), Boolean, String)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Button,System.Action)","name":"Setup(Button, Action)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_Setup_UnityEngine_UIElements_Button_System_Action_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Button,System.Action)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup(UnityEngine.UIElements.Button, System.Action)","nameWithType":"VisualElementExtensions.Setup(Button, Action)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor(UnityEngine.UIElements.VisualElement,System.String,System.String,System.Action{UnityEngine.UIElements.VisualElement})","name":"FindAncestor(VisualElement, String, String, Action<VisualElement>)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_FindAncestor_UnityEngine_UIElements_VisualElement_System_String_System_String_System_Action_UnityEngine_UIElements_VisualElement__","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor(UnityEngine.UIElements.VisualElement,System.String,System.String,System.Action{UnityEngine.UIElements.VisualElement})","name.vb":"FindAncestor(VisualElement, String, String, Action(Of VisualElement))","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor(UnityEngine.UIElements.VisualElement, System.String, System.String, System.Action<UnityEngine.UIElements.VisualElement>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor(UnityEngine.UIElements.VisualElement, System.String, System.String, System.Action(Of UnityEngine.UIElements.VisualElement))","nameWithType":"VisualElementExtensions.FindAncestor(VisualElement, String, String, Action<VisualElement>)","nameWithType.vb":"VisualElementExtensions.FindAncestor(VisualElement, String, String, Action(Of VisualElement))"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot(UnityEngine.UIElements.VisualElement)","name":"GetRoot(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_GetRoot_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot(UnityEngine.UIElements.VisualElement)","nameWithType":"VisualElementExtensions.GetRoot(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor*","name":"DefaultBackgroundColor","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_DefaultBackgroundColor_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.DefaultBackgroundColor","nameWithType":"VisualElementExtensions.DefaultBackgroundColor"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt*","name":"SetEnabledExt","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_SetEnabledExt_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetEnabledExt","nameWithType":"VisualElementExtensions.SetEnabledExt"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt*","name":"SetValueWithoutNotifyExt","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_SetValueWithoutNotifyExt_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.SetValueWithoutNotifyExt","nameWithType":"VisualElementExtensions.SetValueWithoutNotifyExt"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup*","name":"Setup","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_Setup_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.Setup","nameWithType":"VisualElementExtensions.Setup"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor*","name":"FindAncestor","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_FindAncestor_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.FindAncestor","nameWithType":"VisualElementExtensions.FindAncestor"},{"uid":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot*","name":"GetRoot","href":"~/api/AdvancedSceneManager.Editor.Utility.VisualElementExtensions.yml#AdvancedSceneManager_Editor_Utility_VisualElementExtensions_GetRoot_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.VisualElementExtensions.GetRoot","nameWithType":"VisualElementExtensions.GetRoot"}],"api/AdvancedSceneManager.Editor.Utility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility","name":"AdvancedSceneManager.Editor.Utility","href":"~/api/AdvancedSceneManager.Editor.Utility.yml","commentId":"N:AdvancedSceneManager.Editor.Utility","fullName":"AdvancedSceneManager.Editor.Utility","nameWithType":"AdvancedSceneManager.Editor.Utility"}],"api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml":[{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails","name":"CoroutineDiagHelper.SubroutineDetails","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml","commentId":"T:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails","nameWithType":"CoroutineDiagHelper.SubroutineDetails"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.subroutine","name":"subroutine","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_subroutine","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.subroutine","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.subroutine","nameWithType":"CoroutineDiagHelper.SubroutineDetails.subroutine"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.level","name":"level","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_level","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.level","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.level","nameWithType":"CoroutineDiagHelper.SubroutineDetails.level"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.type","name":"type","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_type","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.type","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.type","nameWithType":"CoroutineDiagHelper.SubroutineDetails.type"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isMethod","name":"isMethod","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isMethod","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isMethod","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isMethod","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isMethod"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isValueType","name":"isValueType","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isValueType","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isValueType","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isValueType","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isValueType"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstruction","name":"isDefaultYieldInstruction","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isDefaultYieldInstruction","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstruction","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstruction","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstruction"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstructionComponent","name":"isDefaultYieldInstructionComponent","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isDefaultYieldInstructionComponent","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstructionComponent","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstructionComponent","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isDefaultYieldInstructionComponent"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startTime","name":"startTime","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_startTime","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startTime","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startTime","nameWithType":"CoroutineDiagHelper.SubroutineDetails.startTime"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endTime","name":"endTime","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_endTime","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endTime","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endTime","nameWithType":"CoroutineDiagHelper.SubroutineDetails.endTime"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startFrame","name":"startFrame","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_startFrame","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startFrame","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.startFrame","nameWithType":"CoroutineDiagHelper.SubroutineDetails.startFrame"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endFrame","name":"endFrame","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_endFrame","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endFrame","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.endFrame","nameWithType":"CoroutineDiagHelper.SubroutineDetails.endFrame"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper","name":"helper","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_helper","commentId":"P:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper","nameWithType":"CoroutineDiagHelper.SubroutineDetails.helper"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull","name":"isNull","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isNull","commentId":"P:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isNull"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End","name":"End()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_End","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End()","nameWithType":"CoroutineDiagHelper.SubroutineDetails.End()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_ToString","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString()","nameWithType":"CoroutineDiagHelper.SubroutineDetails.ToString()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.#ctor(System.Object,System.Int32,AdvancedSceneManager.Callbacks.CoroutineDiagHelper,AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","name":"SubroutineDetails(Object, Int32, CoroutineDiagHelper, CoroutineDiagHelper.SubroutineDetails)","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails__ctor_System_Object_System_Int32_AdvancedSceneManager_Callbacks_CoroutineDiagHelper_AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.#ctor(System.Object,System.Int32,AdvancedSceneManager.Callbacks.CoroutineDiagHelper,AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.SubroutineDetails(System.Object, System.Int32, AdvancedSceneManager.Callbacks.CoroutineDiagHelper, AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","nameWithType":"CoroutineDiagHelper.SubroutineDetails.SubroutineDetails(Object, Int32, CoroutineDiagHelper, CoroutineDiagHelper.SubroutineDetails)"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper*","name":"helper","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_helper_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.helper","nameWithType":"CoroutineDiagHelper.SubroutineDetails.helper"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull*","name":"isNull","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_isNull_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.isNull","nameWithType":"CoroutineDiagHelper.SubroutineDetails.isNull"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End*","name":"End","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_End_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.End","nameWithType":"CoroutineDiagHelper.SubroutineDetails.End"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_ToString_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.ToString","nameWithType":"CoroutineDiagHelper.SubroutineDetails.ToString"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.#ctor*","name":"SubroutineDetails","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails__ctor_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails.SubroutineDetails","nameWithType":"CoroutineDiagHelper.SubroutineDetails.SubroutineDetails"}],"api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml":[{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime","name":"SerializableDateTime","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml","commentId":"T:AdvancedSceneManager.Callbacks.SerializableDateTime","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime","nameWithType":"SerializableDateTime"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.Convert(System.DateTime)","name":"Convert(DateTime)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_Convert_System_DateTime_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableDateTime.Convert(System.DateTime)","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.Convert(System.DateTime)","nameWithType":"SerializableDateTime.Convert(DateTime)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack(System.Int64)","name":"ConvertBack(Int64)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_ConvertBack_System_Int64_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack(System.Int64)","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack(System.Int64)","nameWithType":"SerializableDateTime.ConvertBack(Int64)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit(System.DateTime)~AdvancedSceneManager.Callbacks.SerializableDateTime","name":"Implicit(DateTime to SerializableDateTime)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_op_Implicit_System_DateTime__AdvancedSceneManager_Callbacks_SerializableDateTime","commentId":"M:AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit(System.DateTime)~AdvancedSceneManager.Callbacks.SerializableDateTime","name.vb":"Widening(DateTime to SerializableDateTime)","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.Implicit(System.DateTime to AdvancedSceneManager.Callbacks.SerializableDateTime)","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableDateTime.Widening(System.DateTime to AdvancedSceneManager.Callbacks.SerializableDateTime)","nameWithType":"SerializableDateTime.Implicit(DateTime to SerializableDateTime)","nameWithType.vb":"SerializableDateTime.Widening(DateTime to SerializableDateTime)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit(AdvancedSceneManager.Callbacks.SerializableDateTime)~System.DateTime","name":"Implicit(SerializableDateTime to DateTime)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_op_Implicit_AdvancedSceneManager_Callbacks_SerializableDateTime__System_DateTime","commentId":"M:AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit(AdvancedSceneManager.Callbacks.SerializableDateTime)~System.DateTime","name.vb":"Widening(SerializableDateTime to DateTime)","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.Implicit(AdvancedSceneManager.Callbacks.SerializableDateTime to System.DateTime)","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableDateTime.Widening(AdvancedSceneManager.Callbacks.SerializableDateTime to System.DateTime)","nameWithType":"SerializableDateTime.Implicit(SerializableDateTime to DateTime)","nameWithType.vb":"SerializableDateTime.Widening(SerializableDateTime to DateTime)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.ToString(System.String)","name":"ToString(String)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_ToString_System_String_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableDateTime.ToString(System.String)","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.ToString(System.String)","nameWithType":"SerializableDateTime.ToString(String)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.Convert*","name":"Convert","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_Convert_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableDateTime.Convert","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.Convert","nameWithType":"SerializableDateTime.Convert"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack*","name":"ConvertBack","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_ConvertBack_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.ConvertBack","nameWithType":"SerializableDateTime.ConvertBack"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableDateTime.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.Implicit","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableDateTime.Widening","nameWithType":"SerializableDateTime.Implicit","nameWithType.vb":"SerializableDateTime.Widening"},{"uid":"AdvancedSceneManager.Callbacks.SerializableDateTime.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Callbacks.SerializableDateTime.yml#AdvancedSceneManager_Callbacks_SerializableDateTime_ToString_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableDateTime.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableDateTime.ToString","nameWithType":"SerializableDateTime.ToString"}],"api/AdvancedSceneManager.Core.Actions.CallbackAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction","name":"CallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.CallbackAction","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction","nameWithType":"CallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress","nameWithType":"CallbackAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.#ctor(System.Action)","name":"CallbackAction(Action)","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction__ctor_System_Action_","commentId":"M:AdvancedSceneManager.Core.Actions.CallbackAction.#ctor(System.Action)","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.CallbackAction(System.Action)","nameWithType":"CallbackAction.CallbackAction(Action)"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.#ctor(System.Func{System.Collections.IEnumerator})","name":"CallbackAction(Func<IEnumerator>)","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction__ctor_System_Func_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Core.Actions.CallbackAction.#ctor(System.Func{System.Collections.IEnumerator})","name.vb":"CallbackAction(Func(Of IEnumerator))","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.CallbackAction(System.Func<System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Core.Actions.CallbackAction.CallbackAction(System.Func(Of System.Collections.IEnumerator))","nameWithType":"CallbackAction.CallbackAction(Func<IEnumerator>)","nameWithType.vb":"CallbackAction.CallbackAction(Func(Of IEnumerator))"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.CallbackAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"CallbackAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit(System.Action)~AdvancedSceneManager.Core.Actions.CallbackAction","name":"Implicit(Action to CallbackAction)","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_op_Implicit_System_Action__AdvancedSceneManager_Core_Actions_CallbackAction","commentId":"M:AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit(System.Action)~AdvancedSceneManager.Core.Actions.CallbackAction","name.vb":"Widening(Action to CallbackAction)","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.Implicit(System.Action to AdvancedSceneManager.Core.Actions.CallbackAction)","fullName.vb":"AdvancedSceneManager.Core.Actions.CallbackAction.Widening(System.Action to AdvancedSceneManager.Core.Actions.CallbackAction)","nameWithType":"CallbackAction.Implicit(Action to CallbackAction)","nameWithType.vb":"CallbackAction.Widening(Action to CallbackAction)"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit(System.Func{System.Collections.IEnumerator})~AdvancedSceneManager.Core.Actions.CallbackAction","name":"Implicit(Func<IEnumerator> to CallbackAction)","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_op_Implicit_System_Func_System_Collections_IEnumerator___AdvancedSceneManager_Core_Actions_CallbackAction","commentId":"M:AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit(System.Func{System.Collections.IEnumerator})~AdvancedSceneManager.Core.Actions.CallbackAction","name.vb":"Widening(Func(Of IEnumerator) to CallbackAction)","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.Implicit(System.Func<System.Collections.IEnumerator> to AdvancedSceneManager.Core.Actions.CallbackAction)","fullName.vb":"AdvancedSceneManager.Core.Actions.CallbackAction.Widening(System.Func(Of System.Collections.IEnumerator) to AdvancedSceneManager.Core.Actions.CallbackAction)","nameWithType":"CallbackAction.Implicit(Func<IEnumerator> to CallbackAction)","nameWithType.vb":"CallbackAction.Widening(Func(Of IEnumerator) to CallbackAction)"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.reportsProgress","nameWithType":"CallbackAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.#ctor*","name":"CallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CallbackAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.CallbackAction","nameWithType":"CallbackAction.CallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CallbackAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.DoAction","nameWithType":"CallbackAction.DoAction"},{"uid":"AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Core.Actions.CallbackAction.yml#AdvancedSceneManager_Core_Actions_CallbackAction_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CallbackAction.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Core.Actions.CallbackAction.Implicit","fullName.vb":"AdvancedSceneManager.Core.Actions.CallbackAction.Widening","nameWithType":"CallbackAction.Implicit","nameWithType.vb":"CallbackAction.Widening"}],"api/AdvancedSceneManager.Core.Actions.QuickStartupAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.QuickStartupAction","name":"QuickStartupAction","href":"~/api/AdvancedSceneManager.Core.Actions.QuickStartupAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.QuickStartupAction","fullName":"AdvancedSceneManager.Core.Actions.QuickStartupAction","nameWithType":"QuickStartupAction"},{"uid":"AdvancedSceneManager.Core.Actions.QuickStartupAction.#ctor","name":"QuickStartupAction()","href":"~/api/AdvancedSceneManager.Core.Actions.QuickStartupAction.yml#AdvancedSceneManager_Core_Actions_QuickStartupAction__ctor","commentId":"M:AdvancedSceneManager.Core.Actions.QuickStartupAction.#ctor","fullName":"AdvancedSceneManager.Core.Actions.QuickStartupAction.QuickStartupAction()","nameWithType":"QuickStartupAction.QuickStartupAction()"},{"uid":"AdvancedSceneManager.Core.Actions.QuickStartupAction.#ctor*","name":"QuickStartupAction","href":"~/api/AdvancedSceneManager.Core.Actions.QuickStartupAction.yml#AdvancedSceneManager_Core_Actions_QuickStartupAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuickStartupAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuickStartupAction.QuickStartupAction","nameWithType":"QuickStartupAction.QuickStartupAction"}],"api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction","name":"SceneFinishLoadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction","nameWithType":"SceneFinishLoadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","name":"SceneFinishLoadAction(OpenSceneInfo, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction__ctor_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.SceneFinishLoadAction(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneFinishLoadAction.SceneFinishLoadAction(OpenSceneInfo, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name":"SceneFinishLoadAction(Func<OpenSceneInfo>, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction__ctor_System_Func_AdvancedSceneManager_Core_OpenSceneInfo__AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name.vb":"SceneFinishLoadAction(Func(Of OpenSceneInfo), SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.SceneFinishLoadAction(System.Func<AdvancedSceneManager.Core.OpenSceneInfo>, AdvancedSceneManager.Models.SceneCollection)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.SceneFinishLoadAction(System.Func(Of AdvancedSceneManager.Core.OpenSceneInfo), AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneFinishLoadAction.SceneFinishLoadAction(Func<OpenSceneInfo>, SceneCollection)","nameWithType.vb":"SceneFinishLoadAction.SceneFinishLoadAction(Func(Of OpenSceneInfo), SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction(ByRef System.Boolean)","nameWithType":"SceneFinishLoadAction.BeforeDoAction(out Boolean)","nameWithType.vb":"SceneFinishLoadAction.BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneFinishLoadAction.DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor*","name":"SceneFinishLoadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.SceneFinishLoadAction","nameWithType":"SceneFinishLoadAction.SceneFinishLoadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.BeforeDoAction","nameWithType":"SceneFinishLoadAction.BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.yml#AdvancedSceneManager_Core_Actions_SceneFinishLoadAction_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneFinishLoadAction.DoNonOverridenAction","nameWithType":"SceneFinishLoadAction.DoNonOverridenAction"}],"api/AdvancedSceneManager.Core.Actions.StartupAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.StartupAction","name":"StartupAction","href":"~/api/AdvancedSceneManager.Core.Actions.StartupAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.StartupAction","fullName":"AdvancedSceneManager.Core.Actions.StartupAction","nameWithType":"StartupAction"},{"uid":"AdvancedSceneManager.Core.Actions.StartupAction.#ctor(System.Boolean,System.Nullable{UnityEngine.Color},System.Single,System.Single,AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"StartupAction(Boolean, Nullable<Color>, Single, Single, SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.StartupAction.yml#AdvancedSceneManager_Core_Actions_StartupAction__ctor_System_Boolean_System_Nullable_UnityEngine_Color__System_Single_System_Single_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Actions.StartupAction.#ctor(System.Boolean,System.Nullable{UnityEngine.Color},System.Single,System.Single,AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name.vb":"StartupAction(Boolean, Nullable(Of Color), Single, Single, SceneCollection, Boolean)","fullName":"AdvancedSceneManager.Core.Actions.StartupAction.StartupAction(System.Boolean, System.Nullable<UnityEngine.Color>, System.Single, System.Single, AdvancedSceneManager.Models.SceneCollection, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.StartupAction.StartupAction(System.Boolean, System.Nullable(Of UnityEngine.Color), System.Single, System.Single, AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"StartupAction.StartupAction(Boolean, Nullable<Color>, Single, Single, SceneCollection, Boolean)","nameWithType.vb":"StartupAction.StartupAction(Boolean, Nullable(Of Color), Single, Single, SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.StartupAction.#ctor*","name":"StartupAction","href":"~/api/AdvancedSceneManager.Core.Actions.StartupAction.yml#AdvancedSceneManager_Core_Actions_StartupAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.StartupAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.StartupAction.StartupAction","nameWithType":"StartupAction.StartupAction"}],"api/AdvancedSceneManager.Core.Callback.When.yml":[{"uid":"AdvancedSceneManager.Core.Callback.When","name":"Callback.When","href":"~/api/AdvancedSceneManager.Core.Callback.When.yml","commentId":"T:AdvancedSceneManager.Core.Callback.When","fullName":"AdvancedSceneManager.Core.Callback.When","nameWithType":"Callback.When"},{"uid":"AdvancedSceneManager.Core.Callback.When.Before","name":"Before","href":"~/api/AdvancedSceneManager.Core.Callback.When.yml#AdvancedSceneManager_Core_Callback_When_Before","commentId":"F:AdvancedSceneManager.Core.Callback.When.Before","fullName":"AdvancedSceneManager.Core.Callback.When.Before","nameWithType":"Callback.When.Before"},{"uid":"AdvancedSceneManager.Core.Callback.When.After","name":"After","href":"~/api/AdvancedSceneManager.Core.Callback.When.yml#AdvancedSceneManager_Core_Callback_When_After","commentId":"F:AdvancedSceneManager.Core.Callback.When.After","fullName":"AdvancedSceneManager.Core.Callback.When.After","nameWithType":"Callback.When.After"}],"api/AdvancedSceneManager.Core.OpenSceneInfo.yml":[{"uid":"AdvancedSceneManager.Core.OpenSceneInfo","name":"OpenSceneInfo","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml","commentId":"T:AdvancedSceneManager.Core.OpenSceneInfo","fullName":"AdvancedSceneManager.Core.OpenSceneInfo","nameWithType":"OpenSceneInfo"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.scene","name":"scene","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_scene","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.scene","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.scene","nameWithType":"OpenSceneInfo.scene"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.unityScene","name":"unityScene","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_unityScene","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.unityScene","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.unityScene","nameWithType":"OpenSceneInfo.unityScene"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded","name":"isPreloaded","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isPreloaded","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded","nameWithType":"OpenSceneInfo.isPreloaded"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isPersistent","name":"isPersistent","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isPersistent","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isPersistent","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isPersistent","nameWithType":"OpenSceneInfo.isPersistent"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isCollection","name":"isCollection","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isCollection","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isCollection","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isCollection","nameWithType":"OpenSceneInfo.isCollection"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isStandalone","name":"isStandalone","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isStandalone","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isStandalone","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isStandalone","nameWithType":"OpenSceneInfo.isStandalone"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isSpecial","name":"isSpecial","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isSpecial","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isSpecial","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isSpecial","nameWithType":"OpenSceneInfo.isSpecial"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isActive","name":"isActive","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isActive","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isActive","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isActive","nameWithType":"OpenSceneInfo.isActive"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isOpen","name":"isOpen","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isOpen","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.isOpen","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isOpen","nameWithType":"OpenSceneInfo.isOpen"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.sceneManager","name":"sceneManager","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_sceneManager","commentId":"P:AdvancedSceneManager.Core.OpenSceneInfo.sceneManager","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.sceneManager","nameWithType":"OpenSceneInfo.sceneManager"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Object)","name":"Equals(Object)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_System_Object_","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Object)","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Object)","nameWithType":"OpenSceneInfo.Equals(Object)"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode","name":"GetHashCode()","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_GetHashCode","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode()","nameWithType":"OpenSceneInfo.GetHashCode()"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Equals(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"OpenSceneInfo.Equals(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Models.Scene)","name":"Equals(Scene)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(AdvancedSceneManager.Models.Scene)","nameWithType":"OpenSceneInfo.Equals(Scene)"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEngine.SceneManagement.Scene)","name":"Equals(Scene)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEngine.SceneManagement.Scene)","nameWithType":"OpenSceneInfo.Equals(Scene)"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Nullable{UnityEngine.SceneManagement.Scene})","name":"Equals(Nullable<Scene>)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_System_Nullable_UnityEngine_SceneManagement_Scene__","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Nullable{UnityEngine.SceneManagement.Scene})","name.vb":"Equals(Nullable(Of Scene))","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Nullable<UnityEngine.SceneManagement.Scene>)","fullName.vb":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(System.Nullable(Of UnityEngine.SceneManagement.Scene))","nameWithType":"OpenSceneInfo.Equals(Nullable<Scene>)","nameWithType.vb":"OpenSceneInfo.Equals(Nullable(Of Scene))"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEditor.SceneAsset)","name":"Equals(SceneAsset)","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_UnityEditor_SceneAsset_","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEditor.SceneAsset)","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals(UnityEditor.SceneAsset)","nameWithType":"OpenSceneInfo.Equals(SceneAsset)"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_ToString","commentId":"M:AdvancedSceneManager.Core.OpenSceneInfo.ToString","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.ToString()","nameWithType":"OpenSceneInfo.ToString()"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.scene*","name":"scene","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_scene_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.scene","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.scene","nameWithType":"OpenSceneInfo.scene"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.unityScene*","name":"unityScene","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_unityScene_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.unityScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.unityScene","nameWithType":"OpenSceneInfo.unityScene"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded*","name":"isPreloaded","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isPreloaded_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isPreloaded","nameWithType":"OpenSceneInfo.isPreloaded"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isPersistent*","name":"isPersistent","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isPersistent_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isPersistent","nameWithType":"OpenSceneInfo.isPersistent"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isCollection*","name":"isCollection","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isCollection_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isCollection","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isCollection","nameWithType":"OpenSceneInfo.isCollection"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isStandalone*","name":"isStandalone","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isStandalone_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isStandalone","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isStandalone","nameWithType":"OpenSceneInfo.isStandalone"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isSpecial*","name":"isSpecial","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isSpecial_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isSpecial","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isSpecial","nameWithType":"OpenSceneInfo.isSpecial"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isActive*","name":"isActive","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isActive_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isActive","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isActive","nameWithType":"OpenSceneInfo.isActive"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.isOpen*","name":"isOpen","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_isOpen_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.isOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.isOpen","nameWithType":"OpenSceneInfo.isOpen"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.sceneManager*","name":"sceneManager","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_sceneManager_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.sceneManager","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.sceneManager","nameWithType":"OpenSceneInfo.sceneManager"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.Equals*","name":"Equals","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_Equals_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.Equals","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.Equals","nameWithType":"OpenSceneInfo.Equals"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode*","name":"GetHashCode","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_GetHashCode_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.GetHashCode","nameWithType":"OpenSceneInfo.GetHashCode"},{"uid":"AdvancedSceneManager.Core.OpenSceneInfo.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Core.OpenSceneInfo.yml#AdvancedSceneManager_Core_OpenSceneInfo_ToString_","commentId":"Overload:AdvancedSceneManager.Core.OpenSceneInfo.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Core.OpenSceneInfo.ToString","nameWithType":"OpenSceneInfo.ToString"}],"api/AdvancedSceneManager.Core.Phase.yml":[{"uid":"AdvancedSceneManager.Core.Phase","name":"Phase","href":"~/api/AdvancedSceneManager.Core.Phase.yml","commentId":"T:AdvancedSceneManager.Core.Phase","fullName":"AdvancedSceneManager.Core.Phase","nameWithType":"Phase"},{"uid":"AdvancedSceneManager.Core.Phase.CloseCallbacks","name":"CloseCallbacks","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_CloseCallbacks","commentId":"F:AdvancedSceneManager.Core.Phase.CloseCallbacks","fullName":"AdvancedSceneManager.Core.Phase.CloseCallbacks","nameWithType":"Phase.CloseCallbacks"},{"uid":"AdvancedSceneManager.Core.Phase.UnloadScenes","name":"UnloadScenes","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_UnloadScenes","commentId":"F:AdvancedSceneManager.Core.Phase.UnloadScenes","fullName":"AdvancedSceneManager.Core.Phase.UnloadScenes","nameWithType":"Phase.UnloadScenes"},{"uid":"AdvancedSceneManager.Core.Phase.LoadScenes","name":"LoadScenes","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_LoadScenes","commentId":"F:AdvancedSceneManager.Core.Phase.LoadScenes","fullName":"AdvancedSceneManager.Core.Phase.LoadScenes","nameWithType":"Phase.LoadScenes"},{"uid":"AdvancedSceneManager.Core.Phase.OpenCallbacks","name":"OpenCallbacks","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_OpenCallbacks","commentId":"F:AdvancedSceneManager.Core.Phase.OpenCallbacks","fullName":"AdvancedSceneManager.Core.Phase.OpenCallbacks","nameWithType":"Phase.OpenCallbacks"},{"uid":"AdvancedSceneManager.Core.Phase.FinishLoad","name":"FinishLoad","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_FinishLoad","commentId":"F:AdvancedSceneManager.Core.Phase.FinishLoad","fullName":"AdvancedSceneManager.Core.Phase.FinishLoad","nameWithType":"Phase.FinishLoad"},{"uid":"AdvancedSceneManager.Core.Phase.CustomActions","name":"CustomActions","href":"~/api/AdvancedSceneManager.Core.Phase.yml#AdvancedSceneManager_Core_Phase_CustomActions","commentId":"F:AdvancedSceneManager.Core.Phase.CustomActions","fullName":"AdvancedSceneManager.Core.Phase.CustomActions","nameWithType":"Phase.CustomActions"}],"api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen","name":"DefaultLoadingScreen","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.DefaultLoadingScreen","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen","nameWithType":"DefaultLoadingScreen"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.group","name":"group","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_group","commentId":"F:AdvancedSceneManager.Defaults.DefaultLoadingScreen.group","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.group","nameWithType":"DefaultLoadingScreen.group"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.image","name":"image","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_image","commentId":"F:AdvancedSceneManager.Defaults.DefaultLoadingScreen.image","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.image","nameWithType":"DefaultLoadingScreen.image"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.slider","name":"slider","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_slider","commentId":"F:AdvancedSceneManager.Defaults.DefaultLoadingScreen.slider","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.slider","nameWithType":"DefaultLoadingScreen.slider"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.duration","name":"duration","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_duration","commentId":"F:AdvancedSceneManager.Defaults.DefaultLoadingScreen.duration","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.duration","nameWithType":"DefaultLoadingScreen.duration"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.color","name":"color","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_color","commentId":"F:AdvancedSceneManager.Defaults.DefaultLoadingScreen.color","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.color","nameWithType":"DefaultLoadingScreen.color"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"DefaultLoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"DefaultLoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnOpen","nameWithType":"DefaultLoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Defaults.DefaultLoadingScreen.yml#AdvancedSceneManager_Defaults_DefaultLoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.DefaultLoadingScreen.OnClose","nameWithType":"DefaultLoadingScreen.OnClose"}],"api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen","name":"DefaultSplashScreen","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.DefaultSplashScreen","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen","nameWithType":"DefaultSplashScreen"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.group","name":"group","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_group","commentId":"F:AdvancedSceneManager.Defaults.DefaultSplashScreen.group","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.group","nameWithType":"DefaultSplashScreen.group"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.image","name":"image","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_image","commentId":"F:AdvancedSceneManager.Defaults.DefaultSplashScreen.image","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.image","nameWithType":"DefaultSplashScreen.image"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.fadeDuration","name":"fadeDuration","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_fadeDuration","commentId":"F:AdvancedSceneManager.Defaults.DefaultSplashScreen.fadeDuration","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.fadeDuration","nameWithType":"DefaultSplashScreen.fadeDuration"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.waitDuration","name":"waitDuration","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_waitDuration","commentId":"F:AdvancedSceneManager.Defaults.DefaultSplashScreen.waitDuration","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.waitDuration","nameWithType":"DefaultSplashScreen.waitDuration"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen","name":"DisplaySplashScreen()","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_DisplaySplashScreen","commentId":"M:AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen()","nameWithType":"DefaultSplashScreen.DisplaySplashScreen()"},{"uid":"AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen*","name":"DisplaySplashScreen","href":"~/api/AdvancedSceneManager.Defaults.DefaultSplashScreen.yml#AdvancedSceneManager_Defaults_DefaultSplashScreen_DisplaySplashScreen_","commentId":"Overload:AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.DefaultSplashScreen.DisplaySplashScreen","nameWithType":"DefaultSplashScreen.DisplaySplashScreen"}],"api/AdvancedSceneManager.Defaults.yml":[{"uid":"AdvancedSceneManager.Defaults","name":"AdvancedSceneManager.Defaults","href":"~/api/AdvancedSceneManager.Defaults.yml","commentId":"N:AdvancedSceneManager.Defaults","fullName":"AdvancedSceneManager.Defaults","nameWithType":"AdvancedSceneManager.Defaults"}],"api/AdvancedSceneManager.Editor.EditCollectionPopup.yml":[{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup","name":"EditCollectionPopup","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml","commentId":"T:AdvancedSceneManager.Editor.EditCollectionPopup","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup","nameWithType":"EditCollectionPopup"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_path","commentId":"P:AdvancedSceneManager.Editor.EditCollectionPopup.path","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.path","nameWithType":"EditCollectionPopup.path"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.Refresh(AdvancedSceneManager.Models.SceneCollection,System.Action{System.String},System.Action)","name":"Refresh(SceneCollection, Action<String>, Action)","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_Refresh_AdvancedSceneManager_Models_SceneCollection_System_Action_System_String__System_Action_","commentId":"M:AdvancedSceneManager.Editor.EditCollectionPopup.Refresh(AdvancedSceneManager.Models.SceneCollection,System.Action{System.String},System.Action)","name.vb":"Refresh(SceneCollection, Action(Of String), Action)","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.Refresh(AdvancedSceneManager.Models.SceneCollection, System.Action<System.String>, System.Action)","fullName.vb":"AdvancedSceneManager.Editor.EditCollectionPopup.Refresh(AdvancedSceneManager.Models.SceneCollection, System.Action(Of System.String), System.Action)","nameWithType":"EditCollectionPopup.Refresh(SceneCollection, Action<String>, Action)","nameWithType.vb":"EditCollectionPopup.Refresh(SceneCollection, Action(Of String), Action)"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen(AdvancedSceneManager.Editor.EditCollectionPopup)","name":"OnReopen(EditCollectionPopup)","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_OnReopen_AdvancedSceneManager_Editor_EditCollectionPopup_","commentId":"M:AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen(AdvancedSceneManager.Editor.EditCollectionPopup)","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen(AdvancedSceneManager.Editor.EditCollectionPopup)","nameWithType":"EditCollectionPopup.OnReopen(EditCollectionPopup)"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_path_","commentId":"Overload:AdvancedSceneManager.Editor.EditCollectionPopup.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.path","nameWithType":"EditCollectionPopup.path"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.Refresh*","name":"Refresh","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_Refresh_","commentId":"Overload:AdvancedSceneManager.Editor.EditCollectionPopup.Refresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.Refresh","nameWithType":"EditCollectionPopup.Refresh"},{"uid":"AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen*","name":"OnReopen","href":"~/api/AdvancedSceneManager.Editor.EditCollectionPopup.yml#AdvancedSceneManager_Editor_EditCollectionPopup_OnReopen_","commentId":"Overload:AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.EditCollectionPopup.OnReopen","nameWithType":"EditCollectionPopup.OnReopen"}],"api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI","name":"HierarchyGUIUtility.HierarchySceneGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI","nameWithType":"HierarchyGUIUtility.HierarchySceneGUI"}],"api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility","name":"HierarchyGUIUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility","nameWithType":"HierarchyGUIUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI,System.Int32)","name":"AddSceneGUI(HierarchyGUIUtility.HierarchySceneGUI, Int32)","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_AddSceneGUI_AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_HierarchySceneGUI_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI,System.Int32)","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI, System.Int32)","nameWithType":"HierarchyGUIUtility.AddSceneGUI(HierarchyGUIUtility.HierarchySceneGUI, Int32)"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI,System.Int32)","name":"AddGameObjectGUI(HierarchyGUIUtility.HierarchyGameObjectGUI, Int32)","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_AddGameObjectGUI_AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_HierarchyGameObjectGUI_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI,System.Int32)","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI, System.Int32)","nameWithType":"HierarchyGUIUtility.AddGameObjectGUI(HierarchyGUIUtility.HierarchyGameObjectGUI, Int32)"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI)","name":"RemoveSceneGUI(HierarchyGUIUtility.HierarchySceneGUI)","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_RemoveSceneGUI_AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_HierarchySceneGUI_","commentId":"M:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI)","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchySceneGUI)","nameWithType":"HierarchyGUIUtility.RemoveSceneGUI(HierarchyGUIUtility.HierarchySceneGUI)"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI)","name":"RemoveGameObjectGUI(HierarchyGUIUtility.HierarchyGameObjectGUI)","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_RemoveGameObjectGUI_AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_HierarchyGameObjectGUI_","commentId":"M:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI)","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI(AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI)","nameWithType":"HierarchyGUIUtility.RemoveGameObjectGUI(HierarchyGUIUtility.HierarchyGameObjectGUI)"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle","name":"defaultStyle","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_defaultStyle","commentId":"P:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle","nameWithType":"HierarchyGUIUtility.defaultStyle"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint","name":"Repaint()","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_Repaint","commentId":"M:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint()","nameWithType":"HierarchyGUIUtility.Repaint()"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI*","name":"AddSceneGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_AddSceneGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddSceneGUI","nameWithType":"HierarchyGUIUtility.AddSceneGUI"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI*","name":"AddGameObjectGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_AddGameObjectGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.AddGameObjectGUI","nameWithType":"HierarchyGUIUtility.AddGameObjectGUI"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI*","name":"RemoveSceneGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_RemoveSceneGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveSceneGUI","nameWithType":"HierarchyGUIUtility.RemoveSceneGUI"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI*","name":"RemoveGameObjectGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_RemoveGameObjectGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.RemoveGameObjectGUI","nameWithType":"HierarchyGUIUtility.RemoveGameObjectGUI"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle*","name":"defaultStyle","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_defaultStyle_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.defaultStyle","nameWithType":"HierarchyGUIUtility.defaultStyle"},{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint*","name":"Repaint","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.yml#AdvancedSceneManager_Editor_Utility_HierarchyGUIUtility_Repaint_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.Repaint","nameWithType":"HierarchyGUIUtility.Repaint"}],"api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab","name":"SettingsTab","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.SettingsTab","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab","nameWithType":"SettingsTab"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.instance","name":"instance","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_instance","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab.instance","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.instance","nameWithType":"SettingsTab.instance"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.#ctor","name":"SettingsTab()","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__ctor","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.#ctor","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.SettingsTab()","nameWithType":"SettingsTab.SettingsTab()"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder(System.String,System.Int32)","name":"SetHeaderOrder(String, Int32)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_SetHeaderOrder_System_String_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder(System.String,System.Int32)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder(System.String, System.Int32)","nameWithType":"SettingsTab.SetHeaderOrder(String, Int32)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder(System.String)","name":"GetHeaderOrder(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_GetHeaderOrder_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder(System.String)","nameWithType":"SettingsTab.GetHeaderOrder(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent(UnityEngine.UIElements.VisualElement,System.String)","name":"AddHeaderContent(VisualElement, String)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_AddHeaderContent_UnityEngine_UIElements_VisualElement_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent(UnityEngine.UIElements.VisualElement,System.String)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent(UnityEngine.UIElements.VisualElement, System.String)","nameWithType":"SettingsTab.AddHeaderContent(VisualElement, String)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent(UnityEngine.UIElements.VisualElement)","name":"RemoveHeaderContent(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_RemoveHeaderContent_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent(UnityEngine.UIElements.VisualElement)","nameWithType":"SettingsTab.RemoveHeaderContent(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders","name":"DefaultHeaders","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_DefaultHeaders","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders","nameWithType":"SettingsTab.DefaultHeaders"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Add(UnityEngine.UIElements.VisualElement,System.String)","name":"Add(VisualElement, String)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Add_UnityEngine_UIElements_VisualElement_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.Add(UnityEngine.UIElements.VisualElement,System.String)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Add(UnityEngine.UIElements.VisualElement, System.String)","nameWithType":"SettingsTab.Add(VisualElement, String)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer(System.String)","name":"Spacer(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Spacer_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer(System.String)","nameWithType":"SettingsTab.Spacer(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Remove(UnityEngine.UIElements.VisualElement)","name":"Remove(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Remove_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.Utility.SettingsTab.Remove(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Remove(UnityEngine.UIElements.VisualElement)","nameWithType":"SettingsTab.Remove(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.instance*","name":"instance","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_instance_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.instance","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.instance","nameWithType":"SettingsTab.instance"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.#ctor*","name":"SettingsTab","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__ctor_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.SettingsTab","nameWithType":"SettingsTab.SettingsTab"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder*","name":"SetHeaderOrder","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_SetHeaderOrder_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.SetHeaderOrder","nameWithType":"SettingsTab.SetHeaderOrder"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder*","name":"GetHeaderOrder","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_GetHeaderOrder_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.GetHeaderOrder","nameWithType":"SettingsTab.GetHeaderOrder"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent*","name":"AddHeaderContent","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_AddHeaderContent_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.AddHeaderContent","nameWithType":"SettingsTab.AddHeaderContent"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent*","name":"RemoveHeaderContent","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_RemoveHeaderContent_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.RemoveHeaderContent","nameWithType":"SettingsTab.RemoveHeaderContent"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders*","name":"DefaultHeaders","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_DefaultHeaders_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.DefaultHeaders","nameWithType":"SettingsTab.DefaultHeaders"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Add*","name":"Add","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Add_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.Add","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Add","nameWithType":"SettingsTab.Add"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer*","name":"Spacer","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Spacer_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Spacer","nameWithType":"SettingsTab.Spacer"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab.yml#AdvancedSceneManager_Editor_Utility_SettingsTab_Remove_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab.Remove","nameWithType":"SettingsTab.Remove"}],"api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders","name":"SettingsTab._DefaultHeaders","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders","nameWithType":"SettingsTab._DefaultHeaders"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance","name":"Appearance","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance","nameWithType":"SettingsTab._DefaultHeaders.Appearance"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab","name":"Appearance_ScenesTab","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_ScenesTab","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab","nameWithType":"SettingsTab._DefaultHeaders.Appearance_ScenesTab"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader","name":"Appearance_WindowHeader","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_WindowHeader","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader","nameWithType":"SettingsTab._DefaultHeaders.Appearance_WindowHeader"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader","name":"Appearance_CollectionHeader","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_CollectionHeader","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader","nameWithType":"SettingsTab._DefaultHeaders.Appearance_CollectionHeader"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy","name":"Appearance_Hierarchy","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_Hierarchy","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy","nameWithType":"SettingsTab._DefaultHeaders.Appearance_Hierarchy"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options","name":"Options","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options","nameWithType":"SettingsTab._DefaultHeaders.Options"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project","name":"Options_Project","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Project","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project","nameWithType":"SettingsTab._DefaultHeaders.Options_Project"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile","name":"Options_Profile","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Profile","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile","nameWithType":"SettingsTab._DefaultHeaders.Options_Profile"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local","name":"Options_Local","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Local","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local","nameWithType":"SettingsTab._DefaultHeaders.Options_Local"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log","name":"Options_Log","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Log","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log","nameWithType":"SettingsTab._DefaultHeaders.Options_Log"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples","name":"PluginsAndExamples","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins","name":"PluginsAndExamples_Plugins","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Plugins","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments","name":"PluginsAndExamples_Experiments","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Experiments","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples","name":"PluginsAndExamples_Examples","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Examples","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Examples"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist","name":"Blacklist","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Blacklist","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist","nameWithType":"SettingsTab._DefaultHeaders.Blacklist"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections","name":"DynamicCollections","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_DynamicCollections","commentId":"P:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections","nameWithType":"SettingsTab._DefaultHeaders.DynamicCollections"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance*","name":"Appearance","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance","nameWithType":"SettingsTab._DefaultHeaders.Appearance"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab*","name":"Appearance_ScenesTab","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_ScenesTab_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_ScenesTab","nameWithType":"SettingsTab._DefaultHeaders.Appearance_ScenesTab"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader*","name":"Appearance_WindowHeader","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_WindowHeader_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_WindowHeader","nameWithType":"SettingsTab._DefaultHeaders.Appearance_WindowHeader"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader*","name":"Appearance_CollectionHeader","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_CollectionHeader_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_CollectionHeader","nameWithType":"SettingsTab._DefaultHeaders.Appearance_CollectionHeader"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy*","name":"Appearance_Hierarchy","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Appearance_Hierarchy_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Appearance_Hierarchy","nameWithType":"SettingsTab._DefaultHeaders.Appearance_Hierarchy"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options*","name":"Options","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options","nameWithType":"SettingsTab._DefaultHeaders.Options"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project*","name":"Options_Project","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Project_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Project","nameWithType":"SettingsTab._DefaultHeaders.Options_Project"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile*","name":"Options_Profile","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Profile_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Profile","nameWithType":"SettingsTab._DefaultHeaders.Options_Profile"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local*","name":"Options_Local","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Local_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Local","nameWithType":"SettingsTab._DefaultHeaders.Options_Local"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log*","name":"Options_Log","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Options_Log_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Options_Log","nameWithType":"SettingsTab._DefaultHeaders.Options_Log"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples*","name":"PluginsAndExamples","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins*","name":"PluginsAndExamples_Plugins","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Plugins_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Plugins"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments*","name":"PluginsAndExamples_Experiments","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Experiments_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Experiments"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples*","name":"PluginsAndExamples_Examples","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_PluginsAndExamples_Examples_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.PluginsAndExamples_Examples","nameWithType":"SettingsTab._DefaultHeaders.PluginsAndExamples_Examples"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist*","name":"Blacklist","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_Blacklist_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.Blacklist","nameWithType":"SettingsTab._DefaultHeaders.Blacklist"},{"uid":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections*","name":"DynamicCollections","href":"~/api/AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.yml#AdvancedSceneManager_Editor_Utility_SettingsTab__DefaultHeaders_DynamicCollections_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.SettingsTab._DefaultHeaders.DynamicCollections","nameWithType":"SettingsTab._DefaultHeaders.DynamicCollections"}],"api/AdvancedSceneManager.Callbacks.CallbackUtility.yml":[{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility","name":"CallbackUtility","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml","commentId":"T:AdvancedSceneManager.Callbacks.CallbackUtility","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility","nameWithType":"CallbackUtility"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.yieldInstructions","name":"yieldInstructions","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_yieldInstructions","commentId":"F:AdvancedSceneManager.Callbacks.CallbackUtility.yieldInstructions","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.yieldInstructions","nameWithType":"CallbackUtility.yieldInstructions"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.customYieldInstructions","name":"customYieldInstructions","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_customYieldInstructions","commentId":"F:AdvancedSceneManager.Callbacks.CallbackUtility.customYieldInstructions","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.customYieldInstructions","nameWithType":"CallbackUtility.customYieldInstructions"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.delayInstructions","name":"delayInstructions","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_delayInstructions","commentId":"F:AdvancedSceneManager.Callbacks.CallbackUtility.delayInstructions","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.delayInstructions","nameWithType":"CallbackUtility.delayInstructions"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.Open","name":"Open()","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_Open","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.Open","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.Open()","nameWithType":"CallbackUtility.Open()"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.Invoke``1","name":"Invoke<T>()","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_Invoke__1","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.Invoke``1","name.vb":"Invoke(Of T)()","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.Invoke<T>()","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.Invoke(Of T)()","nameWithType":"CallbackUtility.Invoke<T>()","nameWithType.vb":"CallbackUtility.Invoke(Of T)()"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_Open_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.Open","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.Open","nameWithType":"CallbackUtility.Open"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.Invoke*","name":"Invoke","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.yml#AdvancedSceneManager_Callbacks_CallbackUtility_Invoke_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.Invoke","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.Invoke","nameWithType":"CallbackUtility.Invoke"}],"api/AdvancedSceneManager.Callbacks.ICollectionExtraData.yml":[{"uid":"AdvancedSceneManager.Callbacks.ICollectionExtraData","name":"ICollectionExtraData","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionExtraData.yml","commentId":"T:AdvancedSceneManager.Callbacks.ICollectionExtraData","fullName":"AdvancedSceneManager.Callbacks.ICollectionExtraData","nameWithType":"ICollectionExtraData"}],"api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml":[{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan","name":"SerializableTimeSpan","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml","commentId":"T:AdvancedSceneManager.Callbacks.SerializableTimeSpan","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan","nameWithType":"SerializableTimeSpan"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert(System.TimeSpan)","name":"Convert(TimeSpan)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_Convert_System_TimeSpan_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert(System.TimeSpan)","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert(System.TimeSpan)","nameWithType":"SerializableTimeSpan.Convert(TimeSpan)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack(System.Int64)","name":"ConvertBack(Int64)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_ConvertBack_System_Int64_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack(System.Int64)","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack(System.Int64)","nameWithType":"SerializableTimeSpan.ConvertBack(Int64)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit(System.TimeSpan)~AdvancedSceneManager.Callbacks.SerializableTimeSpan","name":"Implicit(TimeSpan to SerializableTimeSpan)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_op_Implicit_System_TimeSpan__AdvancedSceneManager_Callbacks_SerializableTimeSpan","commentId":"M:AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit(System.TimeSpan)~AdvancedSceneManager.Callbacks.SerializableTimeSpan","name.vb":"Widening(TimeSpan to SerializableTimeSpan)","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Implicit(System.TimeSpan to AdvancedSceneManager.Callbacks.SerializableTimeSpan)","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Widening(System.TimeSpan to AdvancedSceneManager.Callbacks.SerializableTimeSpan)","nameWithType":"SerializableTimeSpan.Implicit(TimeSpan to SerializableTimeSpan)","nameWithType.vb":"SerializableTimeSpan.Widening(TimeSpan to SerializableTimeSpan)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit(AdvancedSceneManager.Callbacks.SerializableTimeSpan)~System.TimeSpan","name":"Implicit(SerializableTimeSpan to TimeSpan)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_op_Implicit_AdvancedSceneManager_Callbacks_SerializableTimeSpan__System_TimeSpan","commentId":"M:AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit(AdvancedSceneManager.Callbacks.SerializableTimeSpan)~System.TimeSpan","name.vb":"Widening(SerializableTimeSpan to TimeSpan)","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Implicit(AdvancedSceneManager.Callbacks.SerializableTimeSpan to System.TimeSpan)","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Widening(AdvancedSceneManager.Callbacks.SerializableTimeSpan to System.TimeSpan)","nameWithType":"SerializableTimeSpan.Implicit(SerializableTimeSpan to TimeSpan)","nameWithType.vb":"SerializableTimeSpan.Widening(SerializableTimeSpan to TimeSpan)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString(System.String)","name":"ToString(String)","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_ToString_System_String_","commentId":"M:AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString(System.String)","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString(System.String)","nameWithType":"SerializableTimeSpan.ToString(String)"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert*","name":"Convert","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_Convert_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Convert","nameWithType":"SerializableTimeSpan.Convert"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack*","name":"ConvertBack","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_ConvertBack_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ConvertBack","nameWithType":"SerializableTimeSpan.ConvertBack"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableTimeSpan.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Implicit","fullName.vb":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.Widening","nameWithType":"SerializableTimeSpan.Implicit","nameWithType.vb":"SerializableTimeSpan.Widening"},{"uid":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Callbacks.SerializableTimeSpan.yml#AdvancedSceneManager_Callbacks_SerializableTimeSpan_ToString_","commentId":"Overload:AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.SerializableTimeSpan.ToString","nameWithType":"SerializableTimeSpan.ToString"}],"api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml":[{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1","name":"OpenAndRunCallbackAction<T>","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml","commentId":"T:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1","name.vb":"OpenAndRunCallbackAction(Of T)","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T)","nameWithType":"OpenAndRunCallbackAction<T>","nameWithType.vb":"OpenAndRunCallbackAction(Of T)"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.reportsProgress","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).reportsProgress","nameWithType":"OpenAndRunCallbackAction<T>.reportsProgress","nameWithType.vb":"OpenAndRunCallbackAction(Of T).reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.defaultTimeout","name":"defaultTimeout","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_defaultTimeout","commentId":"F:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.defaultTimeout","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.defaultTimeout","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).defaultTimeout","nameWithType":"OpenAndRunCallbackAction<T>.defaultTimeout","nameWithType.vb":"OpenAndRunCallbackAction(Of T).defaultTimeout"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.#ctor(AdvancedSceneManager.Models.Scene,System.Func{`0,System.Collections.IEnumerator},System.Nullable{System.Single},System.Boolean,System.Action)","name":"OpenAndRunCallbackAction(Scene, Func<T, IEnumerator>, Nullable<Single>, Boolean, Action)","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1__ctor_AdvancedSceneManager_Models_Scene_System_Func__0_System_Collections_IEnumerator__System_Nullable_System_Single__System_Boolean_System_Action_","commentId":"M:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.#ctor(AdvancedSceneManager.Models.Scene,System.Func{`0,System.Collections.IEnumerator},System.Nullable{System.Single},System.Boolean,System.Action)","name.vb":"OpenAndRunCallbackAction(Scene, Func(Of T, IEnumerator), Nullable(Of Single), Boolean, Action)","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.OpenAndRunCallbackAction(AdvancedSceneManager.Models.Scene, System.Func<T, System.Collections.IEnumerator>, System.Nullable<System.Single>, System.Boolean, System.Action)","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).OpenAndRunCallbackAction(AdvancedSceneManager.Models.Scene, System.Func(Of T, System.Collections.IEnumerator), System.Nullable(Of System.Single), System.Boolean, System.Action)","nameWithType":"OpenAndRunCallbackAction<T>.OpenAndRunCallbackAction(Scene, Func<T, IEnumerator>, Nullable<Single>, Boolean, Action)","nameWithType.vb":"OpenAndRunCallbackAction(Of T).OpenAndRunCallbackAction(Scene, Func(Of T, IEnumerator), Nullable(Of Single), Boolean, Action)"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.onMissingCallback","name":"onMissingCallback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_onMissingCallback","commentId":"P:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.onMissingCallback","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.onMissingCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).onMissingCallback","nameWithType":"OpenAndRunCallbackAction<T>.onMissingCallback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).onMissingCallback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.callback","name":"callback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_callback","commentId":"P:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.callback","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.callback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).callback","nameWithType":"OpenAndRunCallbackAction<T>.callback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).callback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.runCallback","name":"runCallback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_runCallback","commentId":"P:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.runCallback","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.runCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).runCallback","nameWithType":"OpenAndRunCallbackAction<T>.runCallback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).runCallback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.isLoadingScreen","name":"isLoadingScreen","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_isLoadingScreen","commentId":"P:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.isLoadingScreen","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.isLoadingScreen","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).isLoadingScreen","nameWithType":"OpenAndRunCallbackAction<T>.isLoadingScreen","nameWithType.vb":"OpenAndRunCallbackAction(Of T).isLoadingScreen"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"OpenAndRunCallbackAction<T>.DoAction(SceneManagerBase)","nameWithType.vb":"OpenAndRunCallbackAction(Of T).DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.reportsProgress","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).reportsProgress","nameWithType":"OpenAndRunCallbackAction<T>.reportsProgress","nameWithType.vb":"OpenAndRunCallbackAction(Of T).reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.#ctor*","name":"OpenAndRunCallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.OpenAndRunCallbackAction","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).OpenAndRunCallbackAction","nameWithType":"OpenAndRunCallbackAction<T>.OpenAndRunCallbackAction","nameWithType.vb":"OpenAndRunCallbackAction(Of T).OpenAndRunCallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.onMissingCallback*","name":"onMissingCallback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_onMissingCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.onMissingCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.onMissingCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).onMissingCallback","nameWithType":"OpenAndRunCallbackAction<T>.onMissingCallback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).onMissingCallback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.callback*","name":"callback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_callback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.callback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.callback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).callback","nameWithType":"OpenAndRunCallbackAction<T>.callback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).callback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.runCallback*","name":"runCallback","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_runCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.runCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.runCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).runCallback","nameWithType":"OpenAndRunCallbackAction<T>.runCallback","nameWithType.vb":"OpenAndRunCallbackAction(Of T).runCallback"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.isLoadingScreen*","name":"isLoadingScreen","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_isLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.isLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.isLoadingScreen","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).isLoadingScreen","nameWithType":"OpenAndRunCallbackAction<T>.isLoadingScreen","nameWithType.vb":"OpenAndRunCallbackAction(Of T).isLoadingScreen"},{"uid":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction-1.yml#AdvancedSceneManager_Core_Actions_OpenAndRunCallbackAction_1_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction`1.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction<T>.DoAction","fullName.vb":"AdvancedSceneManager.Core.Actions.OpenAndRunCallbackAction(Of T).DoAction","nameWithType":"OpenAndRunCallbackAction<T>.DoAction","nameWithType.vb":"OpenAndRunCallbackAction(Of T).DoAction"}],"api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml":[{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1","name":"RunCallbackAndCloseAction<T>","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml","commentId":"T:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1","name.vb":"RunCallbackAndCloseAction(Of T)","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T)","nameWithType":"RunCallbackAndCloseAction<T>","nameWithType.vb":"RunCallbackAndCloseAction(Of T)"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.reportsProgress","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).reportsProgress","nameWithType":"RunCallbackAndCloseAction<T>.reportsProgress","nameWithType.vb":"RunCallbackAndCloseAction(Of T).reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.#ctor(`0,System.Func{`0,System.Collections.IEnumerator},System.Boolean,System.Boolean)","name":"RunCallbackAndCloseAction(T, Func<T, IEnumerator>, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1__ctor__0_System_Func__0_System_Collections_IEnumerator__System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.#ctor(`0,System.Func{`0,System.Collections.IEnumerator},System.Boolean,System.Boolean)","name.vb":"RunCallbackAndCloseAction(T, Func(Of T, IEnumerator), Boolean, Boolean)","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.RunCallbackAndCloseAction(T, System.Func<T, System.Collections.IEnumerator>, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).RunCallbackAndCloseAction(T, System.Func(Of T, System.Collections.IEnumerator), System.Boolean, System.Boolean)","nameWithType":"RunCallbackAndCloseAction<T>.RunCallbackAndCloseAction(T, Func<T, IEnumerator>, Boolean, Boolean)","nameWithType.vb":"RunCallbackAndCloseAction(Of T).RunCallbackAndCloseAction(T, Func(Of T, IEnumerator), Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.closeScene","name":"closeScene","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_closeScene","commentId":"P:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.closeScene","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.closeScene","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).closeScene","nameWithType":"RunCallbackAndCloseAction<T>.closeScene","nameWithType.vb":"RunCallbackAndCloseAction(Of T).closeScene"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.callback","name":"callback","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_callback","commentId":"P:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.callback","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.callback","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).callback","nameWithType":"RunCallbackAndCloseAction<T>.callback","nameWithType.vb":"RunCallbackAndCloseAction(Of T).callback"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.runCallback","name":"runCallback","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_runCallback","commentId":"P:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.runCallback","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.runCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).runCallback","nameWithType":"RunCallbackAndCloseAction<T>.runCallback","nameWithType.vb":"RunCallbackAndCloseAction(Of T).runCallback"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.isLoadingScreen","name":"isLoadingScreen","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_isLoadingScreen","commentId":"P:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.isLoadingScreen","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.isLoadingScreen","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).isLoadingScreen","nameWithType":"RunCallbackAndCloseAction<T>.isLoadingScreen","nameWithType.vb":"RunCallbackAndCloseAction(Of T).isLoadingScreen"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"RunCallbackAndCloseAction<T>.DoAction(SceneManagerBase)","nameWithType.vb":"RunCallbackAndCloseAction(Of T).DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.reportsProgress","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).reportsProgress","nameWithType":"RunCallbackAndCloseAction<T>.reportsProgress","nameWithType.vb":"RunCallbackAndCloseAction(Of T).reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.#ctor*","name":"RunCallbackAndCloseAction","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.RunCallbackAndCloseAction","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).RunCallbackAndCloseAction","nameWithType":"RunCallbackAndCloseAction<T>.RunCallbackAndCloseAction","nameWithType.vb":"RunCallbackAndCloseAction(Of T).RunCallbackAndCloseAction"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.closeScene*","name":"closeScene","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_closeScene_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.closeScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.closeScene","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).closeScene","nameWithType":"RunCallbackAndCloseAction<T>.closeScene","nameWithType.vb":"RunCallbackAndCloseAction(Of T).closeScene"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.callback*","name":"callback","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_callback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.callback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.callback","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).callback","nameWithType":"RunCallbackAndCloseAction<T>.callback","nameWithType.vb":"RunCallbackAndCloseAction(Of T).callback"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.runCallback*","name":"runCallback","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_runCallback_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.runCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.runCallback","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).runCallback","nameWithType":"RunCallbackAndCloseAction<T>.runCallback","nameWithType.vb":"RunCallbackAndCloseAction(Of T).runCallback"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.isLoadingScreen*","name":"isLoadingScreen","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_isLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.isLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.isLoadingScreen","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).isLoadingScreen","nameWithType":"RunCallbackAndCloseAction<T>.isLoadingScreen","nameWithType.vb":"RunCallbackAndCloseAction(Of T).isLoadingScreen"},{"uid":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction-1.yml#AdvancedSceneManager_Core_Actions_RunCallbackAndCloseAction_1_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction`1.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction<T>.DoAction","fullName.vb":"AdvancedSceneManager.Core.Actions.RunCallbackAndCloseAction(Of T).DoAction","nameWithType":"RunCallbackAndCloseAction<T>.DoAction","nameWithType.vb":"RunCallbackAndCloseAction(Of T).DoAction"}],"api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction","name":"SceneUnloadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneUnloadAction","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction","nameWithType":"SceneUnloadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","name":"SceneUnloadAction(OpenSceneInfo, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction__ctor_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.SceneUnloadAction(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneUnloadAction.SceneUnloadAction(OpenSceneInfo, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name":"SceneUnloadAction(Func<OpenSceneInfo>, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction__ctor_System_Func_AdvancedSceneManager_Core_OpenSceneInfo__AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name.vb":"SceneUnloadAction(Func(Of OpenSceneInfo), SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.SceneUnloadAction(System.Func<AdvancedSceneManager.Core.OpenSceneInfo>, AdvancedSceneManager.Models.SceneCollection)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.SceneUnloadAction(System.Func(Of AdvancedSceneManager.Core.OpenSceneInfo), AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneUnloadAction.SceneUnloadAction(Func<OpenSceneInfo>, SceneCollection)","nameWithType.vb":"SceneUnloadAction.SceneUnloadAction(Func(Of OpenSceneInfo), SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction(ByRef System.Boolean)","nameWithType":"SceneUnloadAction.BeforeDoAction(out Boolean)","nameWithType.vb":"SceneUnloadAction.BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneUnloadAction.DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","name":"UnsetPersistentFlag(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_UnsetPersistentFlag_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"SceneUnloadAction.UnsetPersistentFlag(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Core.SceneManagerBase)","name":"Remove(OpenSceneInfo, SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_Remove_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneUnloadAction.Remove(OpenSceneInfo, SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor*","name":"SceneUnloadAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneUnloadAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.SceneUnloadAction","nameWithType":"SceneUnloadAction.SceneUnloadAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.BeforeDoAction","nameWithType":"SceneUnloadAction.BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.DoNonOverridenAction","nameWithType":"SceneUnloadAction.DoNonOverridenAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag*","name":"UnsetPersistentFlag","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_UnsetPersistentFlag_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.UnsetPersistentFlag","nameWithType":"SceneUnloadAction.UnsetPersistentFlag"},{"uid":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Core.Actions.SceneUnloadAction.yml#AdvancedSceneManager_Core_Actions_SceneUnloadAction_Remove_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneUnloadAction.Remove","nameWithType":"SceneUnloadAction.Remove"}],"api/AdvancedSceneManager.Core.Callback.yml":[{"uid":"AdvancedSceneManager.Core.Callback","name":"Callback","href":"~/api/AdvancedSceneManager.Core.Callback.yml","commentId":"T:AdvancedSceneManager.Core.Callback","fullName":"AdvancedSceneManager.Core.Callback","nameWithType":"Callback"},{"uid":"AdvancedSceneManager.Core.Callback.phase","name":"phase","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_phase","commentId":"P:AdvancedSceneManager.Core.Callback.phase","fullName":"AdvancedSceneManager.Core.Callback.phase","nameWithType":"Callback.phase"},{"uid":"AdvancedSceneManager.Core.Callback.when","name":"when","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_when","commentId":"P:AdvancedSceneManager.Core.Callback.when","fullName":"AdvancedSceneManager.Core.Callback.when","nameWithType":"Callback.when"},{"uid":"AdvancedSceneManager.Core.Callback.action","name":"action","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_action","commentId":"P:AdvancedSceneManager.Core.Callback.action","fullName":"AdvancedSceneManager.Core.Callback.action","nameWithType":"Callback.action"},{"uid":"AdvancedSceneManager.Core.Callback.action2","name":"action2","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_action2","commentId":"P:AdvancedSceneManager.Core.Callback.action2","fullName":"AdvancedSceneManager.Core.Callback.action2","nameWithType":"Callback.action2"},{"uid":"AdvancedSceneManager.Core.Callback.enumerator","name":"enumerator","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_enumerator","commentId":"P:AdvancedSceneManager.Core.Callback.enumerator","fullName":"AdvancedSceneManager.Core.Callback.enumerator","nameWithType":"Callback.enumerator"},{"uid":"AdvancedSceneManager.Core.Callback.coroutine","name":"coroutine","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_coroutine","commentId":"P:AdvancedSceneManager.Core.Callback.coroutine","fullName":"AdvancedSceneManager.Core.Callback.coroutine","nameWithType":"Callback.coroutine"},{"uid":"AdvancedSceneManager.Core.Callback.scene","name":"scene","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_scene","commentId":"P:AdvancedSceneManager.Core.Callback.scene","fullName":"AdvancedSceneManager.Core.Callback.scene","nameWithType":"Callback.scene"},{"uid":"AdvancedSceneManager.Core.Callback.op_Implicit(System.Action)~AdvancedSceneManager.Core.Callback","name":"Implicit(Action to Callback)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_op_Implicit_System_Action__AdvancedSceneManager_Core_Callback","commentId":"M:AdvancedSceneManager.Core.Callback.op_Implicit(System.Action)~AdvancedSceneManager.Core.Callback","name.vb":"Widening(Action to Callback)","fullName":"AdvancedSceneManager.Core.Callback.Implicit(System.Action to AdvancedSceneManager.Core.Callback)","fullName.vb":"AdvancedSceneManager.Core.Callback.Widening(System.Action to AdvancedSceneManager.Core.Callback)","nameWithType":"Callback.Implicit(Action to Callback)","nameWithType.vb":"Callback.Widening(Action to Callback)"},{"uid":"AdvancedSceneManager.Core.Callback.op_Implicit(System.Action{AdvancedSceneManager.Core.SceneOperation})~AdvancedSceneManager.Core.Callback","name":"Implicit(Action<SceneOperation> to Callback)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_op_Implicit_System_Action_AdvancedSceneManager_Core_SceneOperation___AdvancedSceneManager_Core_Callback","commentId":"M:AdvancedSceneManager.Core.Callback.op_Implicit(System.Action{AdvancedSceneManager.Core.SceneOperation})~AdvancedSceneManager.Core.Callback","name.vb":"Widening(Action(Of SceneOperation) to Callback)","fullName":"AdvancedSceneManager.Core.Callback.Implicit(System.Action<AdvancedSceneManager.Core.SceneOperation> to AdvancedSceneManager.Core.Callback)","fullName.vb":"AdvancedSceneManager.Core.Callback.Widening(System.Action(Of AdvancedSceneManager.Core.SceneOperation) to AdvancedSceneManager.Core.Callback)","nameWithType":"Callback.Implicit(Action<SceneOperation> to Callback)","nameWithType.vb":"Callback.Widening(Action(Of SceneOperation) to Callback)"},{"uid":"AdvancedSceneManager.Core.Callback.op_Implicit(System.Func{System.Collections.IEnumerator})~AdvancedSceneManager.Core.Callback","name":"Implicit(Func<IEnumerator> to Callback)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_op_Implicit_System_Func_System_Collections_IEnumerator___AdvancedSceneManager_Core_Callback","commentId":"M:AdvancedSceneManager.Core.Callback.op_Implicit(System.Func{System.Collections.IEnumerator})~AdvancedSceneManager.Core.Callback","name.vb":"Widening(Func(Of IEnumerator) to Callback)","fullName":"AdvancedSceneManager.Core.Callback.Implicit(System.Func<System.Collections.IEnumerator> to AdvancedSceneManager.Core.Callback)","fullName.vb":"AdvancedSceneManager.Core.Callback.Widening(System.Func(Of System.Collections.IEnumerator) to AdvancedSceneManager.Core.Callback)","nameWithType":"Callback.Implicit(Func<IEnumerator> to Callback)","nameWithType.vb":"Callback.Widening(Func(Of IEnumerator) to Callback)"},{"uid":"AdvancedSceneManager.Core.Callback.op_Implicit(Lazy.Utility.GlobalCoroutine)~AdvancedSceneManager.Core.Callback","name":"Implicit(GlobalCoroutine to Callback)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_op_Implicit_Lazy_Utility_GlobalCoroutine__AdvancedSceneManager_Core_Callback","commentId":"M:AdvancedSceneManager.Core.Callback.op_Implicit(Lazy.Utility.GlobalCoroutine)~AdvancedSceneManager.Core.Callback","name.vb":"Widening(GlobalCoroutine to Callback)","fullName":"AdvancedSceneManager.Core.Callback.Implicit(Lazy.Utility.GlobalCoroutine to AdvancedSceneManager.Core.Callback)","fullName.vb":"AdvancedSceneManager.Core.Callback.Widening(Lazy.Utility.GlobalCoroutine to AdvancedSceneManager.Core.Callback)","nameWithType":"Callback.Implicit(GlobalCoroutine to Callback)","nameWithType.vb":"Callback.Widening(GlobalCoroutine to Callback)"},{"uid":"AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen","name":"AfterLoadingScreenOpen()","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_AfterLoadingScreenOpen","commentId":"M:AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen","fullName":"AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen()","nameWithType":"Callback.AfterLoadingScreenOpen()"},{"uid":"AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose","name":"BeforeLoadingScreenClose()","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_BeforeLoadingScreenClose","commentId":"M:AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose","fullName":"AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose()","nameWithType":"Callback.BeforeLoadingScreenClose()"},{"uid":"AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Models.Scene)","name":"Before(Phase, Scene)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Before_AdvancedSceneManager_Core_Phase_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase, AdvancedSceneManager.Models.Scene)","nameWithType":"Callback.Before(Phase, Scene)"},{"uid":"AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Models.Scene)","name":"After(Phase, Scene)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_After_AdvancedSceneManager_Core_Phase_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase, AdvancedSceneManager.Models.Scene)","nameWithType":"Callback.After(Phase, Scene)"},{"uid":"AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase)","name":"Before(Phase)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Before_AdvancedSceneManager_Core_Phase_","commentId":"M:AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase)","fullName":"AdvancedSceneManager.Core.Callback.Before(AdvancedSceneManager.Core.Phase)","nameWithType":"Callback.Before(Phase)"},{"uid":"AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase)","name":"After(Phase)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_After_AdvancedSceneManager_Core_Phase_","commentId":"M:AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase)","fullName":"AdvancedSceneManager.Core.Callback.After(AdvancedSceneManager.Core.Phase)","nameWithType":"Callback.After(Phase)"},{"uid":"AdvancedSceneManager.Core.Callback.Do(System.Action)","name":"Do(Action)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_System_Action_","commentId":"M:AdvancedSceneManager.Core.Callback.Do(System.Action)","fullName":"AdvancedSceneManager.Core.Callback.Do(System.Action)","nameWithType":"Callback.Do(Action)"},{"uid":"AdvancedSceneManager.Core.Callback.Do(System.Action{AdvancedSceneManager.Core.SceneOperation})","name":"Do(Action<SceneOperation>)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_System_Action_AdvancedSceneManager_Core_SceneOperation__","commentId":"M:AdvancedSceneManager.Core.Callback.Do(System.Action{AdvancedSceneManager.Core.SceneOperation})","name.vb":"Do(Action(Of SceneOperation))","fullName":"AdvancedSceneManager.Core.Callback.Do(System.Action<AdvancedSceneManager.Core.SceneOperation>)","fullName.vb":"AdvancedSceneManager.Core.Callback.Do(System.Action(Of AdvancedSceneManager.Core.SceneOperation))","nameWithType":"Callback.Do(Action<SceneOperation>)","nameWithType.vb":"Callback.Do(Action(Of SceneOperation))"},{"uid":"AdvancedSceneManager.Core.Callback.Do(System.Func{System.Collections.IEnumerator})","name":"Do(Func<IEnumerator>)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_System_Func_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Core.Callback.Do(System.Func{System.Collections.IEnumerator})","name.vb":"Do(Func(Of IEnumerator))","fullName":"AdvancedSceneManager.Core.Callback.Do(System.Func<System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Core.Callback.Do(System.Func(Of System.Collections.IEnumerator))","nameWithType":"Callback.Do(Func<IEnumerator>)","nameWithType.vb":"Callback.Do(Func(Of IEnumerator))"},{"uid":"AdvancedSceneManager.Core.Callback.Do(Lazy.Utility.GlobalCoroutine)","name":"Do(GlobalCoroutine)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_Lazy_Utility_GlobalCoroutine_","commentId":"M:AdvancedSceneManager.Core.Callback.Do(Lazy.Utility.GlobalCoroutine)","fullName":"AdvancedSceneManager.Core.Callback.Do(Lazy.Utility.GlobalCoroutine)","nameWithType":"Callback.Do(GlobalCoroutine)"},{"uid":"AdvancedSceneManager.Core.Callback.Do(System.Single)","name":"Do(Single)","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_System_Single_","commentId":"M:AdvancedSceneManager.Core.Callback.Do(System.Single)","fullName":"AdvancedSceneManager.Core.Callback.Do(System.Single)","nameWithType":"Callback.Do(Single)"},{"uid":"AdvancedSceneManager.Core.Callback.phase*","name":"phase","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_phase_","commentId":"Overload:AdvancedSceneManager.Core.Callback.phase","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.phase","nameWithType":"Callback.phase"},{"uid":"AdvancedSceneManager.Core.Callback.when*","name":"when","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_when_","commentId":"Overload:AdvancedSceneManager.Core.Callback.when","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.when","nameWithType":"Callback.when"},{"uid":"AdvancedSceneManager.Core.Callback.action*","name":"action","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_action_","commentId":"Overload:AdvancedSceneManager.Core.Callback.action","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.action","nameWithType":"Callback.action"},{"uid":"AdvancedSceneManager.Core.Callback.action2*","name":"action2","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_action2_","commentId":"Overload:AdvancedSceneManager.Core.Callback.action2","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.action2","nameWithType":"Callback.action2"},{"uid":"AdvancedSceneManager.Core.Callback.enumerator*","name":"enumerator","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_enumerator_","commentId":"Overload:AdvancedSceneManager.Core.Callback.enumerator","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.enumerator","nameWithType":"Callback.enumerator"},{"uid":"AdvancedSceneManager.Core.Callback.coroutine*","name":"coroutine","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_coroutine_","commentId":"Overload:AdvancedSceneManager.Core.Callback.coroutine","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.coroutine","nameWithType":"Callback.coroutine"},{"uid":"AdvancedSceneManager.Core.Callback.scene*","name":"scene","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_scene_","commentId":"Overload:AdvancedSceneManager.Core.Callback.scene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.scene","nameWithType":"Callback.scene"},{"uid":"AdvancedSceneManager.Core.Callback.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Core.Callback.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Core.Callback.Implicit","fullName.vb":"AdvancedSceneManager.Core.Callback.Widening","nameWithType":"Callback.Implicit","nameWithType.vb":"Callback.Widening"},{"uid":"AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen*","name":"AfterLoadingScreenOpen","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_AfterLoadingScreenOpen_","commentId":"Overload:AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.AfterLoadingScreenOpen","nameWithType":"Callback.AfterLoadingScreenOpen"},{"uid":"AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose*","name":"BeforeLoadingScreenClose","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_BeforeLoadingScreenClose_","commentId":"Overload:AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.BeforeLoadingScreenClose","nameWithType":"Callback.BeforeLoadingScreenClose"},{"uid":"AdvancedSceneManager.Core.Callback.Before*","name":"Before","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Before_","commentId":"Overload:AdvancedSceneManager.Core.Callback.Before","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.Before","nameWithType":"Callback.Before"},{"uid":"AdvancedSceneManager.Core.Callback.After*","name":"After","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_After_","commentId":"Overload:AdvancedSceneManager.Core.Callback.After","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.After","nameWithType":"Callback.After"},{"uid":"AdvancedSceneManager.Core.Callback.Do*","name":"Do","href":"~/api/AdvancedSceneManager.Core.Callback.yml#AdvancedSceneManager_Core_Callback_Do_","commentId":"Overload:AdvancedSceneManager.Core.Callback.Do","isSpec":"True","fullName":"AdvancedSceneManager.Core.Callback.Do","nameWithType":"Callback.Do"}],"api/AdvancedSceneManager.Core.SceneOperation-1.yml":[{"uid":"AdvancedSceneManager.Core.SceneOperation`1","name":"SceneOperation<ReturnValue>","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml","commentId":"T:AdvancedSceneManager.Core.SceneOperation`1","name.vb":"SceneOperation(Of ReturnValue)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue)","nameWithType":"SceneOperation<ReturnValue>","nameWithType.vb":"SceneOperation(Of ReturnValue)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.done","name":"done","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_done","commentId":"P:AdvancedSceneManager.Core.SceneOperation`1.done","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.done","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).done","nameWithType":"SceneOperation<ReturnValue>.done","nameWithType.vb":"SceneOperation(Of ReturnValue).done"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.value","name":"value","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_value","commentId":"P:AdvancedSceneManager.Core.SceneOperation`1.value","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.value","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).value","nameWithType":"SceneOperation<ReturnValue>.value","nameWithType.vb":"SceneOperation(Of ReturnValue).value"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Return(System.Func{AdvancedSceneManager.Core.SceneOperation{`0},`0})","name":"Return(Func<SceneOperation<ReturnValue>, ReturnValue>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Return_System_Func_AdvancedSceneManager_Core_SceneOperation__0___0__","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Return(System.Func{AdvancedSceneManager.Core.SceneOperation{`0},`0})","name.vb":"Return(Func(Of SceneOperation(Of ReturnValue), ReturnValue))","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Return(System.Func<AdvancedSceneManager.Core.SceneOperation<ReturnValue>, ReturnValue>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Return(System.Func(Of AdvancedSceneManager.Core.SceneOperation(Of ReturnValue), ReturnValue))","nameWithType":"SceneOperation<ReturnValue>.Return(Func<SceneOperation<ReturnValue>, ReturnValue>)","nameWithType.vb":"SceneOperation(Of ReturnValue).Return(Func(Of SceneOperation(Of ReturnValue), ReturnValue))"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithFriendlyText(System.String)","name":"WithFriendlyText(String)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithFriendlyText_System_String_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithFriendlyText(System.String)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithFriendlyText(System.String)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithFriendlyText(System.String)","nameWithType":"SceneOperation<ReturnValue>.WithFriendlyText(String)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithFriendlyText(String)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Open(AdvancedSceneManager.Models.Scene[])","name":"Open(Scene[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Open_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Open(AdvancedSceneManager.Models.Scene[])","name.vb":"Open(Scene())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Open(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Open(AdvancedSceneManager.Models.Scene())","nameWithType":"SceneOperation<ReturnValue>.Open(Scene[])","nameWithType.vb":"SceneOperation(Of ReturnValue).Open(Scene())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Open(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.Boolean)","name":"Open(IEnumerable<Scene>, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Open_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Models_Scene__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Open(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.Boolean)","name.vb":"Open(IEnumerable(Of Scene), Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Open(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Models.Scene>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Open(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Models.Scene), System.Boolean)","nameWithType":"SceneOperation<ReturnValue>.Open(IEnumerable<Scene>, Boolean)","nameWithType.vb":"SceneOperation(Of ReturnValue).Open(IEnumerable(Of Scene), Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Close(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Close_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Close(OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Close(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation<ReturnValue>.Close(OpenSceneInfo[])","nameWithType.vb":"SceneOperation(Of ReturnValue).Close(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Close(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},System.Boolean)","name":"Close(IEnumerable<OpenSceneInfo>, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Close_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Close(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},System.Boolean)","name.vb":"Close(IEnumerable(Of OpenSceneInfo), Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Close(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Close(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo), System.Boolean)","nameWithType":"SceneOperation<ReturnValue>.Close(IEnumerable<OpenSceneInfo>, Boolean)","nameWithType.vb":"SceneOperation(Of ReturnValue).Close(IEnumerable(Of OpenSceneInfo), Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Close(System.Boolean,AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Close(Boolean, OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Close_System_Boolean_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Close(System.Boolean,AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Close(Boolean, OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Close(System.Boolean, AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Close(System.Boolean, AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation<ReturnValue>.Close(Boolean, OpenSceneInfo[])","nameWithType.vb":"SceneOperation(Of ReturnValue).Close(Boolean, OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Reopen(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Reopen_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Reopen(OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Reopen(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation<ReturnValue>.Reopen(OpenSceneInfo[])","nameWithType.vb":"SceneOperation(Of ReturnValue).Reopen(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo})","name":"Reopen(IEnumerable<OpenSceneInfo>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Reopen_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo})","name.vb":"Reopen(IEnumerable(Of OpenSceneInfo))","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Reopen(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Reopen(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo))","nameWithType":"SceneOperation<ReturnValue>.Reopen(IEnumerable<OpenSceneInfo>)","nameWithType.vb":"SceneOperation(Of ReturnValue).Reopen(IEnumerable(Of OpenSceneInfo))"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","name":"WithAction(SceneAction[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithAction_AdvancedSceneManager_Core_Actions_SceneAction___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","name.vb":"WithAction(SceneAction())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithAction(AdvancedSceneManager.Core.Actions.SceneAction())","nameWithType":"SceneOperation<ReturnValue>.WithAction(SceneAction[])","nameWithType.vb":"SceneOperation(Of ReturnValue).WithAction(SceneAction())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithCallback(AdvancedSceneManager.Core.Callback)","name":"WithCallback(Callback)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithCallback_AdvancedSceneManager_Core_Callback_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithCallback(AdvancedSceneManager.Core.Callback)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithCallback(AdvancedSceneManager.Core.Callback)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithCallback(AdvancedSceneManager.Core.Callback)","nameWithType":"SceneOperation<ReturnValue>.WithCallback(Callback)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithCallback(Callback)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithCollection(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"WithCollection(SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithCollection_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithCollection(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithCollection(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithCollection(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"SceneOperation<ReturnValue>.WithCollection(SceneCollection, Boolean)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithCollection(SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen(System.Boolean)","name":"WithLoadingScreen(Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingScreen_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen(System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingScreen(System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingScreen(System.Boolean)","nameWithType":"SceneOperation<ReturnValue>.WithLoadingScreen(Boolean)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingScreen(Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","name":"WithLoadingScreen(Scene)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingScreen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingScreen(AdvancedSceneManager.Models.Scene)","nameWithType":"SceneOperation<ReturnValue>.WithLoadingScreen(Scene)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingScreen(Scene)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithClearUnusedAssets(System.Boolean)","name":"WithClearUnusedAssets(Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithClearUnusedAssets_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithClearUnusedAssets(System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithClearUnusedAssets(System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithClearUnusedAssets(System.Boolean)","nameWithType":"SceneOperation<ReturnValue>.WithClearUnusedAssets(Boolean)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithClearUnusedAssets(Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreenCallback(System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name":"WithLoadingScreenCallback(Action<LoadingScreen>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingScreenCallback_System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreenCallback(System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name.vb":"WithLoadingScreenCallback(Action(Of LoadingScreen))","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingScreenCallback(System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingScreenCallback(System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen))","nameWithType":"SceneOperation<ReturnValue>.WithLoadingScreenCallback(Action<LoadingScreen>)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingScreenCallback(Action(Of LoadingScreen))"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingPriority(UnityEngine.ThreadPriority)","name":"WithLoadingPriority(ThreadPriority)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingPriority_UnityEngine_ThreadPriority_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingPriority(UnityEngine.ThreadPriority)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingPriority(UnityEngine.ThreadPriority)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingPriority(UnityEngine.ThreadPriority)","nameWithType":"SceneOperation<ReturnValue>.WithLoadingPriority(ThreadPriority)","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingPriority(ThreadPriority)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","name":"AsPersistent(SceneCloseBehavior)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_AsPersistent_AdvancedSceneManager_Models_SceneCloseBehavior_","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","nameWithType":"SceneOperation<ReturnValue>.AsPersistent(SceneCloseBehavior)","nameWithType.vb":"SceneOperation(Of ReturnValue).AsPersistent(SceneCloseBehavior)"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Reopen(AdvancedSceneManager.Models.Scene[])","name":"Reopen(Scene[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Reopen_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Reopen(AdvancedSceneManager.Models.Scene[])","name.vb":"Reopen(Scene())","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Reopen(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Reopen(AdvancedSceneManager.Models.Scene())","nameWithType":"SceneOperation<ReturnValue>.Reopen(Scene[])","nameWithType.vb":"SceneOperation(Of ReturnValue).Reopen(Scene())"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene})","name":"Reopen(IEnumerable<Scene>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Reopen_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Models_Scene__","commentId":"M:AdvancedSceneManager.Core.SceneOperation`1.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene})","name.vb":"Reopen(IEnumerable(Of Scene))","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Reopen(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Models.Scene>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Reopen(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Models.Scene))","nameWithType":"SceneOperation<ReturnValue>.Reopen(IEnumerable<Scene>)","nameWithType.vb":"SceneOperation(Of ReturnValue).Reopen(IEnumerable(Of Scene))"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.done*","name":"done","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_done_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.done","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.done","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).done","nameWithType":"SceneOperation<ReturnValue>.done","nameWithType.vb":"SceneOperation(Of ReturnValue).done"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.value*","name":"value","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_value_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.value","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.value","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).value","nameWithType":"SceneOperation<ReturnValue>.value","nameWithType.vb":"SceneOperation(Of ReturnValue).value"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Return*","name":"Return","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Return_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.Return","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Return","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Return","nameWithType":"SceneOperation<ReturnValue>.Return","nameWithType.vb":"SceneOperation(Of ReturnValue).Return"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithFriendlyText*","name":"WithFriendlyText","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithFriendlyText_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithFriendlyText","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithFriendlyText","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithFriendlyText","nameWithType":"SceneOperation<ReturnValue>.WithFriendlyText","nameWithType.vb":"SceneOperation(Of ReturnValue).WithFriendlyText"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Open_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.Open","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Open","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Open","nameWithType":"SceneOperation<ReturnValue>.Open","nameWithType.vb":"SceneOperation(Of ReturnValue).Open"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Close_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.Close","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Close","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Close","nameWithType":"SceneOperation<ReturnValue>.Close","nameWithType.vb":"SceneOperation(Of ReturnValue).Close"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_Reopen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.Reopen","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).Reopen","nameWithType":"SceneOperation<ReturnValue>.Reopen","nameWithType.vb":"SceneOperation(Of ReturnValue).Reopen"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithAction*","name":"WithAction","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithAction_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithAction","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithAction","nameWithType":"SceneOperation<ReturnValue>.WithAction","nameWithType.vb":"SceneOperation(Of ReturnValue).WithAction"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithCallback*","name":"WithCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithCallback","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithCallback","nameWithType":"SceneOperation<ReturnValue>.WithCallback","nameWithType.vb":"SceneOperation(Of ReturnValue).WithCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithCollection*","name":"WithCollection","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithCollection_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithCollection","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithCollection","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithCollection","nameWithType":"SceneOperation<ReturnValue>.WithCollection","nameWithType.vb":"SceneOperation(Of ReturnValue).WithCollection"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen*","name":"WithLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingScreen","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingScreen","nameWithType":"SceneOperation<ReturnValue>.WithLoadingScreen","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithClearUnusedAssets*","name":"WithClearUnusedAssets","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithClearUnusedAssets_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithClearUnusedAssets","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithClearUnusedAssets","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithClearUnusedAssets","nameWithType":"SceneOperation<ReturnValue>.WithClearUnusedAssets","nameWithType.vb":"SceneOperation(Of ReturnValue).WithClearUnusedAssets"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreenCallback*","name":"WithLoadingScreenCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingScreenCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingScreenCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingScreenCallback","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingScreenCallback","nameWithType":"SceneOperation<ReturnValue>.WithLoadingScreenCallback","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingScreenCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.WithLoadingPriority*","name":"WithLoadingPriority","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_WithLoadingPriority_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.WithLoadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.WithLoadingPriority","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).WithLoadingPriority","nameWithType":"SceneOperation<ReturnValue>.WithLoadingPriority","nameWithType.vb":"SceneOperation(Of ReturnValue).WithLoadingPriority"},{"uid":"AdvancedSceneManager.Core.SceneOperation`1.AsPersistent*","name":"AsPersistent","href":"~/api/AdvancedSceneManager.Core.SceneOperation-1.yml#AdvancedSceneManager_Core_SceneOperation_1_AsPersistent_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation`1.AsPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation<ReturnValue>.AsPersistent","fullName.vb":"AdvancedSceneManager.Core.SceneOperation(Of ReturnValue).AsPersistent","nameWithType":"SceneOperation<ReturnValue>.AsPersistent","nameWithType.vb":"SceneOperation(Of ReturnValue).AsPersistent"}],"api/AdvancedSceneManager.Core.StandaloneManager.yml":[{"uid":"AdvancedSceneManager.Core.StandaloneManager","name":"StandaloneManager","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml","commentId":"T:AdvancedSceneManager.Core.StandaloneManager","fullName":"AdvancedSceneManager.Core.StandaloneManager","nameWithType":"StandaloneManager"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.OpenSingle(AdvancedSceneManager.Models.Scene)","name":"OpenSingle(Scene)","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_OpenSingle_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.StandaloneManager.OpenSingle(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.StandaloneManager.OpenSingle(AdvancedSceneManager.Models.Scene)","nameWithType":"StandaloneManager.OpenSingle(Scene)"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.Preload(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"Preload(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_Preload_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.StandaloneManager.Preload(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Core.StandaloneManager.Preload(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"StandaloneManager.Preload(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.preloadedScene","name":"preloadedScene","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_preloadedScene","commentId":"P:AdvancedSceneManager.Core.StandaloneManager.preloadedScene","fullName":"AdvancedSceneManager.Core.StandaloneManager.preloadedScene","nameWithType":"StandaloneManager.preloadedScene"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.OpenSingle*","name":"OpenSingle","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_OpenSingle_","commentId":"Overload:AdvancedSceneManager.Core.StandaloneManager.OpenSingle","isSpec":"True","fullName":"AdvancedSceneManager.Core.StandaloneManager.OpenSingle","nameWithType":"StandaloneManager.OpenSingle"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.Preload*","name":"Preload","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_Preload_","commentId":"Overload:AdvancedSceneManager.Core.StandaloneManager.Preload","isSpec":"True","fullName":"AdvancedSceneManager.Core.StandaloneManager.Preload","nameWithType":"StandaloneManager.Preload"},{"uid":"AdvancedSceneManager.Core.StandaloneManager.preloadedScene*","name":"preloadedScene","href":"~/api/AdvancedSceneManager.Core.StandaloneManager.yml#AdvancedSceneManager_Core_StandaloneManager_preloadedScene_","commentId":"Overload:AdvancedSceneManager.Core.StandaloneManager.preloadedScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.StandaloneManager.preloadedScene","nameWithType":"StandaloneManager.preloadedScene"}],"api/AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChangedHandler.yml":[{"uid":"AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChangedHandler","name":"UtilitySceneManager.ActiveSceneChangedHandler","href":"~/api/AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChangedHandler.yml","commentId":"T:AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChangedHandler","fullName":"AdvancedSceneManager.Core.UtilitySceneManager.ActiveSceneChangedHandler","nameWithType":"UtilitySceneManager.ActiveSceneChangedHandler"}],"api/AdvancedSceneManager.Defaults.Quotes.yml":[{"uid":"AdvancedSceneManager.Defaults.Quotes","name":"Quotes","href":"~/api/AdvancedSceneManager.Defaults.Quotes.yml","commentId":"T:AdvancedSceneManager.Defaults.Quotes","fullName":"AdvancedSceneManager.Defaults.Quotes","nameWithType":"Quotes"},{"uid":"AdvancedSceneManager.Defaults.Quotes.quoteList","name":"quoteList","href":"~/api/AdvancedSceneManager.Defaults.Quotes.yml#AdvancedSceneManager_Defaults_Quotes_quoteList","commentId":"F:AdvancedSceneManager.Defaults.Quotes.quoteList","fullName":"AdvancedSceneManager.Defaults.Quotes.quoteList","nameWithType":"Quotes.quoteList"}],"api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen","name":"VideoLoadingScreen","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.VideoLoadingScreen","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen","nameWithType":"VideoLoadingScreen"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.defaultVideoClip","name":"defaultVideoClip","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_defaultVideoClip","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.defaultVideoClip","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.defaultVideoClip","nameWithType":"VideoLoadingScreen.defaultVideoClip"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.videoClip","name":"videoClip","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_videoClip","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.videoClip","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.videoClip","nameWithType":"VideoLoadingScreen.videoClip"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.group","name":"group","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_group","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.group","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.group","nameWithType":"VideoLoadingScreen.group"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.VideoRenderer","name":"VideoRenderer","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_VideoRenderer","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.VideoRenderer","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.VideoRenderer","nameWithType":"VideoLoadingScreen.VideoRenderer"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.fadeDuration","name":"fadeDuration","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_fadeDuration","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.fadeDuration","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.fadeDuration","nameWithType":"VideoLoadingScreen.fadeDuration"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.videoPlayer","name":"videoPlayer","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_videoPlayer","commentId":"F:AdvancedSceneManager.Defaults.VideoLoadingScreen.videoPlayer","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.videoPlayer","nameWithType":"VideoLoadingScreen.videoPlayer"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"VideoLoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"VideoLoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnOpen","nameWithType":"VideoLoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Defaults.VideoLoadingScreen.yml#AdvancedSceneManager_Defaults_VideoLoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.VideoLoadingScreen.OnClose","nameWithType":"VideoLoadingScreen.OnClose"}],"api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml":[{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits","name":"ObjectField.UxmlTraits","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml","commentId":"T:AdvancedSceneManager.Editor.ObjectField.UxmlTraits","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits","nameWithType":"ObjectField.UxmlTraits"},{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription","name":"uxmlChildElementsDescription","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml#AdvancedSceneManager_Editor_ObjectField_UxmlTraits_uxmlChildElementsDescription","commentId":"P:AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription","nameWithType":"ObjectField.UxmlTraits.uxmlChildElementsDescription"},{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement,UnityEngine.UIElements.IUxmlAttributes,UnityEngine.UIElements.CreationContext)","name":"Init(VisualElement, IUxmlAttributes, CreationContext)","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml#AdvancedSceneManager_Editor_ObjectField_UxmlTraits_Init_UnityEngine_UIElements_VisualElement_UnityEngine_UIElements_IUxmlAttributes_UnityEngine_UIElements_CreationContext_","commentId":"M:AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement,UnityEngine.UIElements.IUxmlAttributes,UnityEngine.UIElements.CreationContext)","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement, UnityEngine.UIElements.IUxmlAttributes, UnityEngine.UIElements.CreationContext)","nameWithType":"ObjectField.UxmlTraits.Init(VisualElement, IUxmlAttributes, CreationContext)"},{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription*","name":"uxmlChildElementsDescription","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml#AdvancedSceneManager_Editor_ObjectField_UxmlTraits_uxmlChildElementsDescription_","commentId":"Overload:AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.uxmlChildElementsDescription","nameWithType":"ObjectField.UxmlTraits.uxmlChildElementsDescription"},{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init*","name":"Init","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlTraits.yml#AdvancedSceneManager_Editor_ObjectField_UxmlTraits_Init_","commentId":"Overload:AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlTraits.Init","nameWithType":"ObjectField.UxmlTraits.Init"}],"api/AdvancedSceneManager.Editor.ObjectField.yml":[{"uid":"AdvancedSceneManager.Editor.ObjectField","name":"ObjectField","href":"~/api/AdvancedSceneManager.Editor.ObjectField.yml","commentId":"T:AdvancedSceneManager.Editor.ObjectField","fullName":"AdvancedSceneManager.Editor.ObjectField","nameWithType":"ObjectField"},{"uid":"AdvancedSceneManager.Editor.ObjectField.isReadOnly","name":"isReadOnly","href":"~/api/AdvancedSceneManager.Editor.ObjectField.yml#AdvancedSceneManager_Editor_ObjectField_isReadOnly","commentId":"P:AdvancedSceneManager.Editor.ObjectField.isReadOnly","fullName":"AdvancedSceneManager.Editor.ObjectField.isReadOnly","nameWithType":"ObjectField.isReadOnly"},{"uid":"AdvancedSceneManager.Editor.ObjectField.#ctor","name":"ObjectField()","href":"~/api/AdvancedSceneManager.Editor.ObjectField.yml#AdvancedSceneManager_Editor_ObjectField__ctor","commentId":"M:AdvancedSceneManager.Editor.ObjectField.#ctor","fullName":"AdvancedSceneManager.Editor.ObjectField.ObjectField()","nameWithType":"ObjectField.ObjectField()"},{"uid":"AdvancedSceneManager.Editor.ObjectField.isReadOnly*","name":"isReadOnly","href":"~/api/AdvancedSceneManager.Editor.ObjectField.yml#AdvancedSceneManager_Editor_ObjectField_isReadOnly_","commentId":"Overload:AdvancedSceneManager.Editor.ObjectField.isReadOnly","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ObjectField.isReadOnly","nameWithType":"ObjectField.isReadOnly"},{"uid":"AdvancedSceneManager.Editor.ObjectField.#ctor*","name":"ObjectField","href":"~/api/AdvancedSceneManager.Editor.ObjectField.yml#AdvancedSceneManager_Editor_ObjectField__ctor_","commentId":"Overload:AdvancedSceneManager.Editor.ObjectField.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ObjectField.ObjectField","nameWithType":"ObjectField.ObjectField"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem","name":"SceneManagerWindow.FooterItem","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem","nameWithType":"SceneManagerWindow.FooterItem"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element","name":"element","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_element","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element","nameWithType":"SceneManagerWindow.FooterItem.element"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left","name":"left","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_left","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left","nameWithType":"SceneManagerWindow.FooterItem.left"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create","name":"Create()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Create","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create()","nameWithType":"SceneManagerWindow.FooterItem.Create()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft","name":"OnLeft()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_OnLeft","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft()","nameWithType":"SceneManagerWindow.FooterItem.OnLeft()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight","name":"OnRight()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_OnRight","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight()","nameWithType":"SceneManagerWindow.FooterItem.OnRight()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button(System.String,System.Action,System.String,System.Action{UnityEngine.UIElements.Button})","name":"Button(String, Action, String, Action<Button>)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Button_System_String_System_Action_System_String_System_Action_UnityEngine_UIElements_Button__","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button(System.String,System.Action,System.String,System.Action{UnityEngine.UIElements.Button})","name.vb":"Button(String, Action, String, Action(Of Button))","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button(System.String, System.Action, System.String, System.Action<UnityEngine.UIElements.Button>)","fullName.vb":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button(System.String, System.Action, System.String, System.Action(Of UnityEngine.UIElements.Button))","nameWithType":"SceneManagerWindow.FooterItem.Button(String, Action, String, Action<Button>)","nameWithType.vb":"SceneManagerWindow.FooterItem.Button(String, Action, String, Action(Of Button))"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element``1(System.String,System.Action{``0},System.String)","name":"Element<T>(String, Action<T>, String)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Element__1_System_String_System_Action___0__System_String_","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element``1(System.String,System.Action{``0},System.String)","name.vb":"Element(Of T)(String, Action(Of T), String)","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element<T>(System.String, System.Action<T>, System.String)","fullName.vb":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element(Of T)(System.String, System.Action(Of T), System.String)","nameWithType":"SceneManagerWindow.FooterItem.Element<T>(String, Action<T>, String)","nameWithType.vb":"SceneManagerWindow.FooterItem.Element(Of T)(String, Action(Of T), String)"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden","name":"Hidden()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Hidden","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden()","nameWithType":"SceneManagerWindow.FooterItem.Hidden()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible(System.Boolean)","name":"Visible(Boolean)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Visible_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible(System.Boolean)","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible(System.Boolean)","nameWithType":"SceneManagerWindow.FooterItem.Visible(Boolean)"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element*","name":"element","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_element_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.element","nameWithType":"SceneManagerWindow.FooterItem.element"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left*","name":"left","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_left_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.left","nameWithType":"SceneManagerWindow.FooterItem.left"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create*","name":"Create","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Create_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Create","nameWithType":"SceneManagerWindow.FooterItem.Create"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft*","name":"OnLeft","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_OnLeft_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnLeft","nameWithType":"SceneManagerWindow.FooterItem.OnLeft"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight*","name":"OnRight","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_OnRight_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.OnRight","nameWithType":"SceneManagerWindow.FooterItem.OnRight"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button*","name":"Button","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Button_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Button","nameWithType":"SceneManagerWindow.FooterItem.Button"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element*","name":"Element","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Element_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Element","nameWithType":"SceneManagerWindow.FooterItem.Element"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden*","name":"Hidden","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Hidden_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Hidden","nameWithType":"SceneManagerWindow.FooterItem.Hidden"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible*","name":"Visible","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.yml#AdvancedSceneManager_Editor_SceneManagerWindow_FooterItem_Visible_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.FooterItem.Visible","nameWithType":"SceneManagerWindow.FooterItem.Visible"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.PostProcess.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.PostProcess","name":"SceneManagerWindow.PostProcess","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.PostProcess.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow.PostProcess","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.PostProcess","nameWithType":"SceneManagerWindow.PostProcess"}],"api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility","name":"BuildEventsUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.BuildEventsUtility","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility","nameWithType":"BuildEventsUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.preBuild","name":"preBuild","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildEventsUtility_preBuild","commentId":"E:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.preBuild","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.preBuild","nameWithType":"BuildEventsUtility.preBuild"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.postBuild","name":"postBuild","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildEventsUtility_postBuild","commentId":"E:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.postBuild","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.postBuild","nameWithType":"BuildEventsUtility.postBuild"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onError","name":"onError","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildEventsUtility_onError","commentId":"E:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onError","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onError","nameWithType":"BuildEventsUtility.onError"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onErrorWithArgs","name":"onErrorWithArgs","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildEventsUtility_onErrorWithArgs","commentId":"E:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onErrorWithArgs","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onErrorWithArgs","nameWithType":"BuildEventsUtility.onErrorWithArgs"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onWarningWithArgs","name":"onWarningWithArgs","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.yml#AdvancedSceneManager_Editor_Utility_BuildEventsUtility_onWarningWithArgs","commentId":"E:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onWarningWithArgs","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.onWarningWithArgs","nameWithType":"BuildEventsUtility.onWarningWithArgs"}],"api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason","name":"BuildSettingsUtility.Reason","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason","nameWithType":"BuildSettingsUtility.Reason"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.None","name":"None","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_Reason_None","commentId":"F:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.None","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.None","nameWithType":"BuildSettingsUtility.Reason.None"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.NotIncludedInProfile","name":"NotIncludedInProfile","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_Reason_NotIncludedInProfile","commentId":"F:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.NotIncludedInProfile","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.NotIncludedInProfile","nameWithType":"BuildSettingsUtility.Reason.NotIncludedInProfile"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IncludedInProfile","name":"IncludedInProfile","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_Reason_IncludedInProfile","commentId":"F:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IncludedInProfile","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IncludedInProfile","nameWithType":"BuildSettingsUtility.Reason.IncludedInProfile"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IsAddressable","name":"IsAddressable","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_Reason_IsAddressable","commentId":"F:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IsAddressable","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.IsAddressable","nameWithType":"BuildSettingsUtility.Reason.IsAddressable"},{"uid":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.Overriden","name":"Overriden","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.yml#AdvancedSceneManager_Editor_Utility_BuildSettingsUtility_Reason_Overriden","commentId":"F:AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.Overriden","fullName":"AdvancedSceneManager.Editor.Utility.BuildSettingsUtility.Reason.Overriden","nameWithType":"BuildSettingsUtility.Reason.Overriden"}],"api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting","name":"PersistentSceneInEditorUtility.OpenInEditorSetting","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save","name":"Save()","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_Save","commentId":"M:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save()","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.Save()"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.name","name":"name","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_name","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.name","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.name","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.name"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.scene","name":"scene","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_scene","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.scene","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.scene","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.scene"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.option","name":"option","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_option","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.option","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.option","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.option"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.list","name":"list","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_list","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.list","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.list","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.list"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save*","name":"Save","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorSetting_Save_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorSetting.Save","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorSetting.Save"}],"api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility","name":"PersistentSceneInEditorUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility","nameWithType":"PersistentSceneInEditorUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption(AdvancedSceneManager.Models.Scene)","name":"GetPersistentOption(Scene)","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_GetPersistentOption_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption(AdvancedSceneManager.Models.Scene)","nameWithType":"PersistentSceneInEditorUtility.GetPersistentOption(Scene)"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"OpenAssociatedPersistentScenes(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenAssociatedPersistentScenes_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes(AdvancedSceneManager.Models.Scene)","name":"GetAssociatedScenes(Scene)","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_GetAssociatedScenes_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes(AdvancedSceneManager.Models.Scene)","nameWithType":"PersistentSceneInEditorUtility.GetAssociatedScenes(Scene)"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent(UnityEngine.SceneManagement.Scene)","name":"IsPersistent(Scene)","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_IsPersistent_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent(UnityEngine.SceneManagement.Scene)","nameWithType":"PersistentSceneInEditorUtility.IsPersistent(Scene)"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption*","name":"GetPersistentOption","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_GetPersistentOption_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetPersistentOption","nameWithType":"PersistentSceneInEditorUtility.GetPersistentOption"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes*","name":"OpenAssociatedPersistentScenes","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenAssociatedPersistentScenes_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes","nameWithType":"PersistentSceneInEditorUtility.OpenAssociatedPersistentScenes"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes*","name":"GetAssociatedScenes","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_GetAssociatedScenes_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.GetAssociatedScenes","nameWithType":"PersistentSceneInEditorUtility.GetAssociatedScenes"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent*","name":"IsPersistent","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_IsPersistent_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.IsPersistent","nameWithType":"PersistentSceneInEditorUtility.IsPersistent"}],"api/AdvancedSceneManager.Models.SceneCloseBehavior.yml":[{"uid":"AdvancedSceneManager.Models.SceneCloseBehavior","name":"SceneCloseBehavior","href":"~/api/AdvancedSceneManager.Models.SceneCloseBehavior.yml","commentId":"T:AdvancedSceneManager.Models.SceneCloseBehavior","fullName":"AdvancedSceneManager.Models.SceneCloseBehavior","nameWithType":"SceneCloseBehavior"},{"uid":"AdvancedSceneManager.Models.SceneCloseBehavior.Close","name":"Close","href":"~/api/AdvancedSceneManager.Models.SceneCloseBehavior.yml#AdvancedSceneManager_Models_SceneCloseBehavior_Close","commentId":"F:AdvancedSceneManager.Models.SceneCloseBehavior.Close","fullName":"AdvancedSceneManager.Models.SceneCloseBehavior.Close","nameWithType":"SceneCloseBehavior.Close"},{"uid":"AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenIfNextCollectionAlsoContainsScene","name":"KeepOpenIfNextCollectionAlsoContainsScene","href":"~/api/AdvancedSceneManager.Models.SceneCloseBehavior.yml#AdvancedSceneManager_Models_SceneCloseBehavior_KeepOpenIfNextCollectionAlsoContainsScene","commentId":"F:AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenIfNextCollectionAlsoContainsScene","fullName":"AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenIfNextCollectionAlsoContainsScene","nameWithType":"SceneCloseBehavior.KeepOpenIfNextCollectionAlsoContainsScene"},{"uid":"AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenAlways","name":"KeepOpenAlways","href":"~/api/AdvancedSceneManager.Models.SceneCloseBehavior.yml#AdvancedSceneManager_Models_SceneCloseBehavior_KeepOpenAlways","commentId":"F:AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenAlways","fullName":"AdvancedSceneManager.Models.SceneCloseBehavior.KeepOpenAlways","nameWithType":"SceneCloseBehavior.KeepOpenAlways"}],"api/AdvancedSceneManager.Models.SceneCollection.yml":[{"uid":"AdvancedSceneManager.Models.SceneCollection","name":"SceneCollection","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml","commentId":"T:AdvancedSceneManager.Models.SceneCollection","fullName":"AdvancedSceneManager.Models.SceneCollection","nameWithType":"SceneCollection"},{"uid":"AdvancedSceneManager.Models.SceneCollection.PropertyChanged","name":"PropertyChanged","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_PropertyChanged","commentId":"E:AdvancedSceneManager.Models.SceneCollection.PropertyChanged","fullName":"AdvancedSceneManager.Models.SceneCollection.PropertyChanged","nameWithType":"SceneCollection.PropertyChanged"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged","name":"OnPropertyChanged()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OnPropertyChanged","commentId":"M:AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged","fullName":"AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged()","nameWithType":"SceneCollection.OnPropertyChanged()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Count","name":"Count","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Count","commentId":"P:AdvancedSceneManager.Models.SceneCollection.Count","fullName":"AdvancedSceneManager.Models.SceneCollection.Count","nameWithType":"SceneCollection.Count"},{"uid":"AdvancedSceneManager.Models.SceneCollection.IsReadOnly","name":"IsReadOnly","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_IsReadOnly","commentId":"P:AdvancedSceneManager.Models.SceneCollection.IsReadOnly","fullName":"AdvancedSceneManager.Models.SceneCollection.IsReadOnly","nameWithType":"SceneCollection.IsReadOnly"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Item(System.Int32)","name":"Item[Int32]","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Item_System_Int32_","commentId":"P:AdvancedSceneManager.Models.SceneCollection.Item(System.Int32)","name.vb":"Item(Int32)","fullName":"AdvancedSceneManager.Models.SceneCollection.Item[System.Int32]","fullName.vb":"AdvancedSceneManager.Models.SceneCollection.Item(System.Int32)","nameWithType":"SceneCollection.Item[Int32]","nameWithType.vb":"SceneCollection.Item(Int32)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Contains(AdvancedSceneManager.Models.Scene)","name":"Contains(Scene)","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Contains_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Contains(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Models.SceneCollection.Contains(AdvancedSceneManager.Models.Scene)","nameWithType":"SceneCollection.Contains(Scene)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.GetEnumerator","name":"GetEnumerator()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_GetEnumerator","commentId":"M:AdvancedSceneManager.Models.SceneCollection.GetEnumerator","fullName":"AdvancedSceneManager.Models.SceneCollection.GetEnumerator()","nameWithType":"SceneCollection.GetEnumerator()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.name","name":"name","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_name","commentId":"P:AdvancedSceneManager.Models.SceneCollection.name","fullName":"AdvancedSceneManager.Models.SceneCollection.name","nameWithType":"SceneCollection.name"},{"uid":"AdvancedSceneManager.Models.SceneCollection.title","name":"title","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_title","commentId":"P:AdvancedSceneManager.Models.SceneCollection.title","fullName":"AdvancedSceneManager.Models.SceneCollection.title","nameWithType":"SceneCollection.title"},{"uid":"AdvancedSceneManager.Models.SceneCollection.extraData","name":"extraData","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_extraData","commentId":"P:AdvancedSceneManager.Models.SceneCollection.extraData","fullName":"AdvancedSceneManager.Models.SceneCollection.extraData","nameWithType":"SceneCollection.extraData"},{"uid":"AdvancedSceneManager.Models.SceneCollection.isIncluded","name":"isIncluded","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_isIncluded","commentId":"P:AdvancedSceneManager.Models.SceneCollection.isIncluded","fullName":"AdvancedSceneManager.Models.SceneCollection.isIncluded","nameWithType":"SceneCollection.isIncluded"},{"uid":"AdvancedSceneManager.Models.SceneCollection.scenes","name":"scenes","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_scenes","commentId":"P:AdvancedSceneManager.Models.SceneCollection.scenes","fullName":"AdvancedSceneManager.Models.SceneCollection.scenes","nameWithType":"SceneCollection.scenes"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingScreen","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingScreen","commentId":"P:AdvancedSceneManager.Models.SceneCollection.loadingScreen","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingScreen","nameWithType":"SceneCollection.loadingScreen"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage","name":"loadingScreenUsage","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingScreenUsage","commentId":"P:AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage","nameWithType":"SceneCollection.loadingScreenUsage"},{"uid":"AdvancedSceneManager.Models.SceneCollection.activeScene","name":"activeScene","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_activeScene","commentId":"P:AdvancedSceneManager.Models.SceneCollection.activeScene","fullName":"AdvancedSceneManager.Models.SceneCollection.activeScene","nameWithType":"SceneCollection.activeScene"},{"uid":"AdvancedSceneManager.Models.SceneCollection.startupOption","name":"startupOption","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_startupOption","commentId":"P:AdvancedSceneManager.Models.SceneCollection.startupOption","fullName":"AdvancedSceneManager.Models.SceneCollection.startupOption","nameWithType":"SceneCollection.startupOption"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingPriority","name":"loadingPriority","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingPriority","commentId":"P:AdvancedSceneManager.Models.SceneCollection.loadingPriority","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingPriority","nameWithType":"SceneCollection.loadingPriority"},{"uid":"AdvancedSceneManager.Models.SceneCollection.hasScenes","name":"hasScenes","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_hasScenes","commentId":"P:AdvancedSceneManager.Models.SceneCollection.hasScenes","fullName":"AdvancedSceneManager.Models.SceneCollection.hasScenes","nameWithType":"SceneCollection.hasScenes"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Tag(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneTag)","name":"Tag(Scene, SceneTag)","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Tag_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneTag_","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Tag(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneTag)","fullName":"AdvancedSceneManager.Models.SceneCollection.Tag(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.SceneTag)","nameWithType":"SceneCollection.Tag(Scene, SceneTag)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Open","name":"Open()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Open","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Open","fullName":"AdvancedSceneManager.Models.SceneCollection.Open()","nameWithType":"SceneCollection.Open()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OpenOrReopen","name":"OpenOrReopen()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OpenOrReopen","commentId":"M:AdvancedSceneManager.Models.SceneCollection.OpenOrReopen","fullName":"AdvancedSceneManager.Models.SceneCollection.OpenOrReopen()","nameWithType":"SceneCollection.OpenOrReopen()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Toggle","name":"Toggle()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Toggle","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Toggle","fullName":"AdvancedSceneManager.Models.SceneCollection.Toggle()","nameWithType":"SceneCollection.Toggle()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Toggle(System.Boolean)","name":"Toggle(Boolean)","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Toggle_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Toggle(System.Boolean)","fullName":"AdvancedSceneManager.Models.SceneCollection.Toggle(System.Boolean)","nameWithType":"SceneCollection.Toggle(Boolean)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Reopen","name":"Reopen()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Reopen","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Reopen","fullName":"AdvancedSceneManager.Models.SceneCollection.Reopen()","nameWithType":"SceneCollection.Reopen()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Close","name":"Close()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Close","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Close","fullName":"AdvancedSceneManager.Models.SceneCollection.Close()","nameWithType":"SceneCollection.Close()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.IsOpen","name":"IsOpen()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_IsOpen","commentId":"M:AdvancedSceneManager.Models.SceneCollection.IsOpen","fullName":"AdvancedSceneManager.Models.SceneCollection.IsOpen()","nameWithType":"SceneCollection.IsOpen()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OpenEvent","name":"OpenEvent()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OpenEvent","commentId":"M:AdvancedSceneManager.Models.SceneCollection.OpenEvent","fullName":"AdvancedSceneManager.Models.SceneCollection.OpenEvent()","nameWithType":"SceneCollection.OpenEvent()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent","name":"ToggleEvent()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ToggleEvent","commentId":"M:AdvancedSceneManager.Models.SceneCollection.ToggleEvent","fullName":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent()","nameWithType":"SceneCollection.ToggleEvent()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent(System.Boolean)","name":"ToggleEvent(Boolean)","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ToggleEvent_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.SceneCollection.ToggleEvent(System.Boolean)","fullName":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent(System.Boolean)","nameWithType":"SceneCollection.ToggleEvent(Boolean)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ReopenEvent","name":"ReopenEvent()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ReopenEvent","commentId":"M:AdvancedSceneManager.Models.SceneCollection.ReopenEvent","fullName":"AdvancedSceneManager.Models.SceneCollection.ReopenEvent()","nameWithType":"SceneCollection.ReopenEvent()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.CloseEvent","name":"CloseEvent()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_CloseEvent","commentId":"M:AdvancedSceneManager.Models.SceneCollection.CloseEvent","fullName":"AdvancedSceneManager.Models.SceneCollection.CloseEvent()","nameWithType":"SceneCollection.CloseEvent()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.AllScenes","name":"AllScenes()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_AllScenes","commentId":"M:AdvancedSceneManager.Models.SceneCollection.AllScenes","fullName":"AdvancedSceneManager.Models.SceneCollection.AllScenes()","nameWithType":"SceneCollection.AllScenes()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.AllScenePaths","name":"AllScenePaths()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_AllScenePaths","commentId":"M:AdvancedSceneManager.Models.SceneCollection.AllScenePaths","fullName":"AdvancedSceneManager.Models.SceneCollection.AllScenePaths()","nameWithType":"SceneCollection.AllScenePaths()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.FindProfile","name":"FindProfile()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_FindProfile","commentId":"M:AdvancedSceneManager.Models.SceneCollection.FindProfile","fullName":"AdvancedSceneManager.Models.SceneCollection.FindProfile()","nameWithType":"SceneCollection.FindProfile()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Find(System.String,System.Boolean)","name":"Find(String, Boolean)","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Find_System_String_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.SceneCollection.Find(System.String,System.Boolean)","fullName":"AdvancedSceneManager.Models.SceneCollection.Find(System.String, System.Boolean)","nameWithType":"SceneCollection.Find(String, Boolean)"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ExtraData``1","name":"ExtraData<T>()","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ExtraData__1","commentId":"M:AdvancedSceneManager.Models.SceneCollection.ExtraData``1","name.vb":"ExtraData(Of T)()","fullName":"AdvancedSceneManager.Models.SceneCollection.ExtraData<T>()","fullName.vb":"AdvancedSceneManager.Models.SceneCollection.ExtraData(Of T)()","nameWithType":"SceneCollection.ExtraData<T>()","nameWithType.vb":"SceneCollection.ExtraData(Of T)()"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged*","name":"OnPropertyChanged","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OnPropertyChanged_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.OnPropertyChanged","nameWithType":"SceneCollection.OnPropertyChanged"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Count*","name":"Count","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Count_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Count","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Count","nameWithType":"SceneCollection.Count"},{"uid":"AdvancedSceneManager.Models.SceneCollection.IsReadOnly*","name":"IsReadOnly","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_IsReadOnly_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.IsReadOnly","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.IsReadOnly","nameWithType":"SceneCollection.IsReadOnly"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Item*","name":"Item","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Item_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Item","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Item","nameWithType":"SceneCollection.Item"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Contains*","name":"Contains","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Contains_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Contains","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Contains","nameWithType":"SceneCollection.Contains"},{"uid":"AdvancedSceneManager.Models.SceneCollection.GetEnumerator*","name":"GetEnumerator","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_GetEnumerator_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.GetEnumerator","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.GetEnumerator","nameWithType":"SceneCollection.GetEnumerator"},{"uid":"AdvancedSceneManager.Models.SceneCollection.name*","name":"name","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_name_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.name","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.name","nameWithType":"SceneCollection.name"},{"uid":"AdvancedSceneManager.Models.SceneCollection.title*","name":"title","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_title_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.title","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.title","nameWithType":"SceneCollection.title"},{"uid":"AdvancedSceneManager.Models.SceneCollection.extraData*","name":"extraData","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_extraData_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.extraData","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.extraData","nameWithType":"SceneCollection.extraData"},{"uid":"AdvancedSceneManager.Models.SceneCollection.isIncluded*","name":"isIncluded","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_isIncluded_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.isIncluded","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.isIncluded","nameWithType":"SceneCollection.isIncluded"},{"uid":"AdvancedSceneManager.Models.SceneCollection.scenes*","name":"scenes","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_scenes_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.scenes","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.scenes","nameWithType":"SceneCollection.scenes"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingScreen*","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingScreen_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.loadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingScreen","nameWithType":"SceneCollection.loadingScreen"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage*","name":"loadingScreenUsage","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingScreenUsage_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingScreenUsage","nameWithType":"SceneCollection.loadingScreenUsage"},{"uid":"AdvancedSceneManager.Models.SceneCollection.activeScene*","name":"activeScene","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_activeScene_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.activeScene","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.activeScene","nameWithType":"SceneCollection.activeScene"},{"uid":"AdvancedSceneManager.Models.SceneCollection.startupOption*","name":"startupOption","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_startupOption_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.startupOption","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.startupOption","nameWithType":"SceneCollection.startupOption"},{"uid":"AdvancedSceneManager.Models.SceneCollection.loadingPriority*","name":"loadingPriority","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_loadingPriority_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.loadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.loadingPriority","nameWithType":"SceneCollection.loadingPriority"},{"uid":"AdvancedSceneManager.Models.SceneCollection.hasScenes*","name":"hasScenes","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_hasScenes_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.hasScenes","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.hasScenes","nameWithType":"SceneCollection.hasScenes"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Tag*","name":"Tag","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Tag_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Tag","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Tag","nameWithType":"SceneCollection.Tag"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Open_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Open","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Open","nameWithType":"SceneCollection.Open"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OpenOrReopen*","name":"OpenOrReopen","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OpenOrReopen_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.OpenOrReopen","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.OpenOrReopen","nameWithType":"SceneCollection.OpenOrReopen"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Toggle_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Toggle","nameWithType":"SceneCollection.Toggle"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Reopen_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Reopen","nameWithType":"SceneCollection.Reopen"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Close_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Close","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Close","nameWithType":"SceneCollection.Close"},{"uid":"AdvancedSceneManager.Models.SceneCollection.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_IsOpen_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.IsOpen","nameWithType":"SceneCollection.IsOpen"},{"uid":"AdvancedSceneManager.Models.SceneCollection.OpenEvent*","name":"OpenEvent","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_OpenEvent_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.OpenEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.OpenEvent","nameWithType":"SceneCollection.OpenEvent"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent*","name":"ToggleEvent","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ToggleEvent_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.ToggleEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.ToggleEvent","nameWithType":"SceneCollection.ToggleEvent"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ReopenEvent*","name":"ReopenEvent","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ReopenEvent_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.ReopenEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.ReopenEvent","nameWithType":"SceneCollection.ReopenEvent"},{"uid":"AdvancedSceneManager.Models.SceneCollection.CloseEvent*","name":"CloseEvent","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_CloseEvent_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.CloseEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.CloseEvent","nameWithType":"SceneCollection.CloseEvent"},{"uid":"AdvancedSceneManager.Models.SceneCollection.AllScenes*","name":"AllScenes","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_AllScenes_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.AllScenes","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.AllScenes","nameWithType":"SceneCollection.AllScenes"},{"uid":"AdvancedSceneManager.Models.SceneCollection.AllScenePaths*","name":"AllScenePaths","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_AllScenePaths_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.AllScenePaths","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.AllScenePaths","nameWithType":"SceneCollection.AllScenePaths"},{"uid":"AdvancedSceneManager.Models.SceneCollection.FindProfile*","name":"FindProfile","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_FindProfile_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.FindProfile","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.FindProfile","nameWithType":"SceneCollection.FindProfile"},{"uid":"AdvancedSceneManager.Models.SceneCollection.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_Find_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.Find","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.Find","nameWithType":"SceneCollection.Find"},{"uid":"AdvancedSceneManager.Models.SceneCollection.ExtraData*","name":"ExtraData","href":"~/api/AdvancedSceneManager.Models.SceneCollection.yml#AdvancedSceneManager_Models_SceneCollection_ExtraData_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollection.ExtraData","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollection.ExtraData","nameWithType":"SceneCollection.ExtraData"}],"api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml":[{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility","name":"CanvasSortOrderUtility","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml","commentId":"T:AdvancedSceneManager.Utility.CanvasSortOrderUtility","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility","nameWithType":"CanvasSortOrderUtility"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove(UnityEngine.Canvas)","name":"Remove(Canvas)","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_Remove_UnityEngine_Canvas_","commentId":"M:AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove(UnityEngine.Canvas)","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove(UnityEngine.Canvas)","nameWithType":"CanvasSortOrderUtility.Remove(Canvas)"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop(UnityEngine.Canvas)","name":"PutOnTop(Canvas)","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_PutOnTop_UnityEngine_Canvas_","commentId":"M:AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop(UnityEngine.Canvas)","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop(UnityEngine.Canvas)","nameWithType":"CanvasSortOrderUtility.PutOnTop(Canvas)"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom(UnityEngine.Canvas)","name":"PutAtBottom(Canvas)","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_PutAtBottom_UnityEngine_Canvas_","commentId":"M:AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom(UnityEngine.Canvas)","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom(UnityEngine.Canvas)","nameWithType":"CanvasSortOrderUtility.PutAtBottom(Canvas)"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure(UnityEngine.Canvas,UnityEngine.Canvas,UnityEngine.Canvas)","name":"MakeSure(Canvas, Canvas, Canvas)","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_MakeSure_UnityEngine_Canvas_UnityEngine_Canvas_UnityEngine_Canvas_","commentId":"M:AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure(UnityEngine.Canvas,UnityEngine.Canvas,UnityEngine.Canvas)","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure(UnityEngine.Canvas, UnityEngine.Canvas, UnityEngine.Canvas)","nameWithType":"CanvasSortOrderUtility.MakeSure(Canvas, Canvas, Canvas)"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_Remove_","commentId":"Overload:AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.Remove","nameWithType":"CanvasSortOrderUtility.Remove"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop*","name":"PutOnTop","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_PutOnTop_","commentId":"Overload:AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop","isSpec":"True","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutOnTop","nameWithType":"CanvasSortOrderUtility.PutOnTop"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom*","name":"PutAtBottom","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_PutAtBottom_","commentId":"Overload:AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom","isSpec":"True","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.PutAtBottom","nameWithType":"CanvasSortOrderUtility.PutAtBottom"},{"uid":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure*","name":"MakeSure","href":"~/api/AdvancedSceneManager.Utility.CanvasSortOrderUtility.yml#AdvancedSceneManager_Utility_CanvasSortOrderUtility_MakeSure_","commentId":"Overload:AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure","isSpec":"True","fullName":"AdvancedSceneManager.Utility.CanvasSortOrderUtility.MakeSure","nameWithType":"CanvasSortOrderUtility.MakeSure"}],"api/AdvancedSceneManager.Utility.DefaultSceneUtility.yml":[{"uid":"AdvancedSceneManager.Utility.DefaultSceneUtility","name":"DefaultSceneUtility","href":"~/api/AdvancedSceneManager.Utility.DefaultSceneUtility.yml","commentId":"T:AdvancedSceneManager.Utility.DefaultSceneUtility","fullName":"AdvancedSceneManager.Utility.DefaultSceneUtility","nameWithType":"DefaultSceneUtility"},{"uid":"AdvancedSceneManager.Utility.DefaultSceneUtility.Name","name":"Name","href":"~/api/AdvancedSceneManager.Utility.DefaultSceneUtility.yml#AdvancedSceneManager_Utility_DefaultSceneUtility_Name","commentId":"F:AdvancedSceneManager.Utility.DefaultSceneUtility.Name","fullName":"AdvancedSceneManager.Utility.DefaultSceneUtility.Name","nameWithType":"DefaultSceneUtility.Name"},{"uid":"AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene(UnityEngine.SceneManagement.Scene)","name":"IsDefaultScene(Scene)","href":"~/api/AdvancedSceneManager.Utility.DefaultSceneUtility.yml#AdvancedSceneManager_Utility_DefaultSceneUtility_IsDefaultScene_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene(UnityEngine.SceneManagement.Scene)","nameWithType":"DefaultSceneUtility.IsDefaultScene(Scene)"},{"uid":"AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene*","name":"IsDefaultScene","href":"~/api/AdvancedSceneManager.Utility.DefaultSceneUtility.yml#AdvancedSceneManager_Utility_DefaultSceneUtility_IsDefaultScene_","commentId":"Overload:AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DefaultSceneUtility.IsDefaultScene","nameWithType":"DefaultSceneUtility.IsDefaultScene"}],"api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml":[{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility","name":"SceneCollectionUtility","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml","commentId":"T:AdvancedSceneManager.Utility.SceneCollectionUtility","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility","nameWithType":"SceneCollectionUtility"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Create(System.String,AdvancedSceneManager.Models.Profile)","name":"Create(String, Profile)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Create_System_String_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Create(System.String,AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Create(System.String, AdvancedSceneManager.Models.Profile)","nameWithType":"SceneCollectionUtility.Create(String, Profile)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Remove(AdvancedSceneManager.Models.SceneCollection)","name":"Remove(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Remove_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Remove(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Remove(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCollectionUtility.Remove(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes(AdvancedSceneManager.Models.SceneCollection)","name":"RemoveNullScenes(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_RemoveNullScenes_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCollectionUtility.RemoveNullScenes(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.String)","name":"Find(IEnumerable<Scene>, String)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Find_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Models_Scene__System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.String)","name.vb":"Find(IEnumerable(Of Scene), String)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Models.Scene>, System.String)","fullName.vb":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Models.Scene), System.String)","nameWithType":"SceneCollectionUtility.Find(IEnumerable<Scene>, String)","nameWithType.vb":"SceneCollectionUtility.Find(IEnumerable(Of Scene), String)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{UnityEngine.SceneManagement.Scene},System.String)","name":"Find(IEnumerable<Scene>, String)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Find_System_Collections_Generic_IEnumerable_UnityEngine_SceneManagement_Scene__System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{UnityEngine.SceneManagement.Scene},System.String)","name.vb":"Find(IEnumerable(Of Scene), String)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable<UnityEngine.SceneManagement.Scene>, System.String)","fullName.vb":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable(Of UnityEngine.SceneManagement.Scene), System.String)","nameWithType":"SceneCollectionUtility.Find(IEnumerable<Scene>, String)","nameWithType.vb":"SceneCollectionUtility.Find(IEnumerable(Of Scene), String)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.Scene)","name":"Find(IEnumerable<OpenSceneInfo>, Scene)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Find_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.Scene)","name.vb":"Find(IEnumerable(Of OpenSceneInfo), Scene)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>, AdvancedSceneManager.Models.Scene)","fullName.vb":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo), AdvancedSceneManager.Models.Scene)","nameWithType":"SceneCollectionUtility.Find(IEnumerable<OpenSceneInfo>, Scene)","nameWithType.vb":"SceneCollectionUtility.Find(IEnumerable(Of OpenSceneInfo), Scene)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},UnityEngine.SceneManagement.Scene)","name":"Find(IEnumerable<OpenSceneInfo>, Scene)","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Find_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},UnityEngine.SceneManagement.Scene)","name.vb":"Find(IEnumerable(Of OpenSceneInfo), Scene)","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>, UnityEngine.SceneManagement.Scene)","fullName.vb":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo), UnityEngine.SceneManagement.Scene)","nameWithType":"SceneCollectionUtility.Find(IEnumerable<OpenSceneInfo>, Scene)","nameWithType.vb":"SceneCollectionUtility.Find(IEnumerable(Of OpenSceneInfo), Scene)"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Create*","name":"Create","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Create_","commentId":"Overload:AdvancedSceneManager.Utility.SceneCollectionUtility.Create","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Create","nameWithType":"SceneCollectionUtility.Create"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Remove_","commentId":"Overload:AdvancedSceneManager.Utility.SceneCollectionUtility.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Remove","nameWithType":"SceneCollectionUtility.Remove"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes*","name":"RemoveNullScenes","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_RemoveNullScenes_","commentId":"Overload:AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.RemoveNullScenes","nameWithType":"SceneCollectionUtility.RemoveNullScenes"},{"uid":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Utility.SceneCollectionUtility.yml#AdvancedSceneManager_Utility_SceneCollectionUtility_Find_","commentId":"Overload:AdvancedSceneManager.Utility.SceneCollectionUtility.Find","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneCollectionUtility.Find","nameWithType":"SceneCollectionUtility.Find"}],"api/AdvancedSceneManager.Utility.SceneDataUtility.yml":[{"uid":"AdvancedSceneManager.Utility.SceneDataUtility","name":"SceneDataUtility","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml","commentId":"T:AdvancedSceneManager.Utility.SceneDataUtility","fullName":"AdvancedSceneManager.Utility.SceneDataUtility","nameWithType":"SceneDataUtility"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Enumerate``1(System.String)","name":"Enumerate<T>(String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Enumerate__1_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Enumerate``1(System.String)","name.vb":"Enumerate(Of T)(String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Enumerate<T>(System.String)","fullName.vb":"AdvancedSceneManager.Utility.SceneDataUtility.Enumerate(Of T)(System.String)","nameWithType":"SceneDataUtility.Enumerate<T>(String)","nameWithType.vb":"SceneDataUtility.Enumerate(Of T)(String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Get``1(AdvancedSceneManager.Models.Scene,System.String,``0)","name":"Get<T>(Scene, String, T)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Get__1_AdvancedSceneManager_Models_Scene_System_String___0_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Get``1(AdvancedSceneManager.Models.Scene,System.String,``0)","name.vb":"Get(Of T)(Scene, String, T)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Get<T>(AdvancedSceneManager.Models.Scene, System.String, T)","fullName.vb":"AdvancedSceneManager.Utility.SceneDataUtility.Get(Of T)(AdvancedSceneManager.Models.Scene, System.String, T)","nameWithType":"SceneDataUtility.Get<T>(Scene, String, T)","nameWithType.vb":"SceneDataUtility.Get(Of T)(Scene, String, T)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(AdvancedSceneManager.Models.Scene,System.String)","name":"GetDirect(Scene, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_GetDirect_AdvancedSceneManager_Models_Scene_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(AdvancedSceneManager.Models.Scene,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(AdvancedSceneManager.Models.Scene, System.String)","nameWithType":"SceneDataUtility.GetDirect(Scene, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Set``1(AdvancedSceneManager.Models.Scene,System.String,``0)","name":"Set<T>(Scene, String, T)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Set__1_AdvancedSceneManager_Models_Scene_System_String___0_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Set``1(AdvancedSceneManager.Models.Scene,System.String,``0)","name.vb":"Set(Of T)(Scene, String, T)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Set<T>(AdvancedSceneManager.Models.Scene, System.String, T)","fullName.vb":"AdvancedSceneManager.Utility.SceneDataUtility.Set(Of T)(AdvancedSceneManager.Models.Scene, System.String, T)","nameWithType":"SceneDataUtility.Set<T>(Scene, String, T)","nameWithType.vb":"SceneDataUtility.Set(Of T)(Scene, String, T)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(AdvancedSceneManager.Models.Scene,System.String,System.String)","name":"SetDirect(Scene, String, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_SetDirect_AdvancedSceneManager_Models_Scene_System_String_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(AdvancedSceneManager.Models.Scene,System.String,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(AdvancedSceneManager.Models.Scene, System.String, System.String)","nameWithType":"SceneDataUtility.SetDirect(Scene, String, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Unset(AdvancedSceneManager.Models.Scene,System.String)","name":"Unset(Scene, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Unset_AdvancedSceneManager_Models_Scene_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Unset(AdvancedSceneManager.Models.Scene,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Unset(AdvancedSceneManager.Models.Scene, System.String)","nameWithType":"SceneDataUtility.Unset(Scene, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Get``1(System.String,System.String,``0)","name":"Get<T>(String, String, T)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Get__1_System_String_System_String___0_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Get``1(System.String,System.String,``0)","name.vb":"Get(Of T)(String, String, T)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Get<T>(System.String, System.String, T)","fullName.vb":"AdvancedSceneManager.Utility.SceneDataUtility.Get(Of T)(System.String, System.String, T)","nameWithType":"SceneDataUtility.Get<T>(String, String, T)","nameWithType.vb":"SceneDataUtility.Get(Of T)(String, String, T)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(System.String,System.String)","name":"GetDirect(String, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_GetDirect_System_String_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(System.String,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect(System.String, System.String)","nameWithType":"SceneDataUtility.GetDirect(String, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Set``1(System.String,System.String,``0)","name":"Set<T>(String, String, T)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Set__1_System_String_System_String___0_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Set``1(System.String,System.String,``0)","name.vb":"Set(Of T)(String, String, T)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Set<T>(System.String, System.String, T)","fullName.vb":"AdvancedSceneManager.Utility.SceneDataUtility.Set(Of T)(System.String, System.String, T)","nameWithType":"SceneDataUtility.Set<T>(String, String, T)","nameWithType.vb":"SceneDataUtility.Set(Of T)(String, String, T)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(System.String,System.String,System.String)","name":"SetDirect(String, String, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_SetDirect_System_String_System_String_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(System.String,System.String,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect(System.String, System.String, System.String)","nameWithType":"SceneDataUtility.SetDirect(String, String, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Unset(System.String,System.String)","name":"Unset(String, String)","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Unset_System_String_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneDataUtility.Unset(System.String,System.String)","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Unset(System.String, System.String)","nameWithType":"SceneDataUtility.Unset(String, String)"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Enumerate*","name":"Enumerate","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Enumerate_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.Enumerate","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Enumerate","nameWithType":"SceneDataUtility.Enumerate"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Get*","name":"Get","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Get_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.Get","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Get","nameWithType":"SceneDataUtility.Get"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect*","name":"GetDirect","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_GetDirect_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.GetDirect","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.GetDirect","nameWithType":"SceneDataUtility.GetDirect"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Set*","name":"Set","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Set_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.Set","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Set","nameWithType":"SceneDataUtility.Set"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect*","name":"SetDirect","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_SetDirect_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.SetDirect","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.SetDirect","nameWithType":"SceneDataUtility.SetDirect"},{"uid":"AdvancedSceneManager.Utility.SceneDataUtility.Unset*","name":"Unset","href":"~/api/AdvancedSceneManager.Utility.SceneDataUtility.yml#AdvancedSceneManager_Utility_SceneDataUtility_Unset_","commentId":"Overload:AdvancedSceneManager.Utility.SceneDataUtility.Unset","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneDataUtility.Unset","nameWithType":"SceneDataUtility.Unset"}],"api/AdvancedSceneManager.Utility.SceneHelper.yml":[{"uid":"AdvancedSceneManager.Utility.SceneHelper","name":"SceneHelper","href":"~/api/AdvancedSceneManager.Utility.SceneHelper.yml","commentId":"T:AdvancedSceneManager.Utility.SceneHelper","fullName":"AdvancedSceneManager.Utility.SceneHelper","nameWithType":"SceneHelper"},{"uid":"AdvancedSceneManager.Utility.SceneHelper.current","name":"current","href":"~/api/AdvancedSceneManager.Utility.SceneHelper.yml#AdvancedSceneManager_Utility_SceneHelper_current","commentId":"P:AdvancedSceneManager.Utility.SceneHelper.current","fullName":"AdvancedSceneManager.Utility.SceneHelper.current","nameWithType":"SceneHelper.current"},{"uid":"AdvancedSceneManager.Utility.SceneHelper.current*","name":"current","href":"~/api/AdvancedSceneManager.Utility.SceneHelper.yml#AdvancedSceneManager_Utility_SceneHelper_current_","commentId":"Overload:AdvancedSceneManager.Utility.SceneHelper.current","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneHelper.current","nameWithType":"SceneHelper.current"}],"api/AdvancedSceneManager.Utility.SceneUtility.yml":[{"uid":"AdvancedSceneManager.Utility.SceneUtility","name":"SceneUtility","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml","commentId":"T:AdvancedSceneManager.Utility.SceneUtility","fullName":"AdvancedSceneManager.Utility.SceneUtility","nameWithType":"SceneUtility"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes","name":"GetAllOpenUnityScenes()","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_GetAllOpenUnityScenes","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes","fullName":"AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes()","nameWithType":"SceneUtility.GetAllOpenUnityScenes()"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.isStartupScene","name":"isStartupScene","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_isStartupScene","commentId":"P:AdvancedSceneManager.Utility.SceneUtility.isStartupScene","fullName":"AdvancedSceneManager.Utility.SceneUtility.isStartupScene","nameWithType":"SceneUtility.isStartupScene"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes","name":"hasAnyScenes","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_hasAnyScenes","commentId":"P:AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes","fullName":"AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes","nameWithType":"SceneUtility.hasAnyScenes"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.sceneCount","name":"sceneCount","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_sceneCount","commentId":"P:AdvancedSceneManager.Utility.SceneUtility.sceneCount","fullName":"AdvancedSceneManager.Utility.SceneUtility.sceneCount","nameWithType":"SceneUtility.sceneCount"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject,AdvancedSceneManager.Core.OpenSceneInfo)","name":"Move(GameObject, OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Move_UnityEngine_GameObject_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject,AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject, AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"SceneUtility.Move(GameObject, OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject,UnityEngine.SceneManagement.Scene)","name":"Move(GameObject, Scene)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Move_UnityEngine_GameObject_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject,UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Move(UnityEngine.GameObject, UnityEngine.SceneManagement.Scene)","nameWithType":"SceneUtility.Move(GameObject, Scene)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.CreateDynamic(System.String,UnityEngine.SceneManagement.LocalPhysicsMode)","name":"CreateDynamic(String, LocalPhysicsMode)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_CreateDynamic_System_String_UnityEngine_SceneManagement_LocalPhysicsMode_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.CreateDynamic(System.String,UnityEngine.SceneManagement.LocalPhysicsMode)","fullName":"AdvancedSceneManager.Utility.SceneUtility.CreateDynamic(System.String, UnityEngine.SceneManagement.LocalPhysicsMode)","nameWithType":"SceneUtility.CreateDynamic(String, LocalPhysicsMode)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder(System.Action{AdvancedSceneManager.Models.Scene},AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean)","name":"CreateInCurrentFolder(Action<Scene>, SceneCollection, Nullable<Int32>, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_CreateInCurrentFolder_System_Action_AdvancedSceneManager_Models_Scene__AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Int32__System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder(System.Action{AdvancedSceneManager.Models.Scene},AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean)","name.vb":"CreateInCurrentFolder(Action(Of Scene), SceneCollection, Nullable(Of Int32), Boolean, Boolean)","fullName":"AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder(System.Action<AdvancedSceneManager.Models.Scene>, AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Int32>, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder(System.Action(Of AdvancedSceneManager.Models.Scene), AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Int32), System.Boolean, System.Boolean)","nameWithType":"SceneUtility.CreateInCurrentFolder(Action<Scene>, SceneCollection, Nullable<Int32>, Boolean, Boolean)","nameWithType.vb":"SceneUtility.CreateInCurrentFolder(Action(Of Scene), SceneCollection, Nullable(Of Int32), Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Create(System.Action{AdvancedSceneManager.Models.Scene},AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean)","name":"Create(Action<Scene>, SceneCollection, Nullable<Int32>, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Create_System_Action_AdvancedSceneManager_Models_Scene__AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Int32__System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Create(System.Action{AdvancedSceneManager.Models.Scene},AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean)","name.vb":"Create(Action(Of Scene), SceneCollection, Nullable(Of Int32), Boolean, Boolean)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Create(System.Action<AdvancedSceneManager.Models.Scene>, AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Int32>, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.Create(System.Action(Of AdvancedSceneManager.Models.Scene), AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Int32), System.Boolean, System.Boolean)","nameWithType":"SceneUtility.Create(Action<Scene>, SceneCollection, Nullable<Int32>, Boolean, Boolean)","nameWithType.vb":"SceneUtility.Create(Action(Of Scene), SceneCollection, Nullable(Of Int32), Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Create(System.String,AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean,System.Boolean)","name":"Create(String, SceneCollection, Nullable<Int32>, Boolean, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Create_System_String_AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Int32__System_Boolean_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Create(System.String,AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32},System.Boolean,System.Boolean,System.Boolean)","name.vb":"Create(String, SceneCollection, Nullable(Of Int32), Boolean, Boolean, Boolean)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Create(System.String, AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Int32>, System.Boolean, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.Create(System.String, AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Int32), System.Boolean, System.Boolean, System.Boolean)","nameWithType":"SceneUtility.Create(String, SceneCollection, Nullable<Int32>, Boolean, Boolean, Boolean)","nameWithType.vb":"SceneUtility.Create(String, SceneCollection, Nullable(Of Int32), Boolean, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Remove(System.String)","name":"Remove(String)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Remove_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Remove(System.String)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Remove(System.String)","nameWithType":"SceneUtility.Remove(String)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Remove(AdvancedSceneManager.Models.Scene)","name":"Remove(Scene)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Remove_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Remove(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Remove(AdvancedSceneManager.Models.Scene)","nameWithType":"SceneUtility.Remove(Scene)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.String)","name":"FindOpen(String)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_FindOpen_System_String_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.String)","fullName":"AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.String)","nameWithType":"SceneUtility.FindOpen(String)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.Func{AdvancedSceneManager.Models.Scene,System.Boolean})","name":"FindOpen(Func<Scene, Boolean>)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_FindOpen_System_Func_AdvancedSceneManager_Models_Scene_System_Boolean__","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.Func{AdvancedSceneManager.Models.Scene,System.Boolean})","name.vb":"FindOpen(Func(Of Scene, Boolean))","fullName":"AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.Func<AdvancedSceneManager.Models.Scene, System.Boolean>)","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.FindOpen(System.Func(Of AdvancedSceneManager.Models.Scene, System.Boolean))","nameWithType":"SceneUtility.FindOpen(Func<Scene, Boolean>)","nameWithType.vb":"SceneUtility.FindOpen(Func(Of Scene, Boolean))"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Find(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name":"Find(String, SceneCollection, Profile)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Find_System_String_AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Find(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Find(System.String, AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","nameWithType":"SceneUtility.Find(String, SceneCollection, Profile)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Find(System.Func{AdvancedSceneManager.Models.Scene,System.Boolean},AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name":"Find(Func<Scene, Boolean>, SceneCollection, Profile)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Find_System_Func_AdvancedSceneManager_Models_Scene_System_Boolean__AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Find(System.Func{AdvancedSceneManager.Models.Scene,System.Boolean},AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name.vb":"Find(Func(Of Scene, Boolean), SceneCollection, Profile)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Find(System.Func<AdvancedSceneManager.Models.Scene, System.Boolean>, AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.Find(System.Func(Of AdvancedSceneManager.Models.Scene, System.Boolean), AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","nameWithType":"SceneUtility.Find(Func<Scene, Boolean>, SceneCollection, Profile)","nameWithType.vb":"SceneUtility.Find(Func(Of Scene, Boolean), SceneCollection, Profile)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene(UnityEngine.GameObject[])","name":"MoveToNewScene(GameObject[])","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_MoveToNewScene_UnityEngine_GameObject___","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene(UnityEngine.GameObject[])","name.vb":"MoveToNewScene(GameObject())","fullName":"AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene(UnityEngine.GameObject[])","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene(UnityEngine.GameObject())","nameWithType":"SceneUtility.MoveToNewScene(GameObject[])","nameWithType.vb":"SceneUtility.MoveToNewScene(GameObject())"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.MergeScenes(System.String[])","name":"MergeScenes(String[])","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_MergeScenes_System_String___","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.MergeScenes(System.String[])","name.vb":"MergeScenes(String())","fullName":"AdvancedSceneManager.Utility.SceneUtility.MergeScenes(System.String[])","fullName.vb":"AdvancedSceneManager.Utility.SceneUtility.MergeScenes(System.String())","nameWithType":"SceneUtility.MergeScenes(String[])","nameWithType.vb":"SceneUtility.MergeScenes(String())"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.GameObject)","name":"Scene(GameObject)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Scene_UnityEngine_GameObject_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.GameObject)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.GameObject)","nameWithType":"SceneUtility.Scene(GameObject)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.Component)","name":"Scene(Component)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Scene_UnityEngine_Component_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.Component)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.Component)","nameWithType":"SceneUtility.Scene(Component)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.SceneManagement.Scene)","name":"Scene(Scene)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Scene_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.SceneUtility.Scene(UnityEngine.SceneManagement.Scene)","nameWithType":"SceneUtility.Scene(Scene)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.FindASMScene(UnityEditor.SceneAsset)","name":"FindASMScene(SceneAsset)","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_FindASMScene_UnityEditor_SceneAsset_","commentId":"M:AdvancedSceneManager.Utility.SceneUtility.FindASMScene(UnityEditor.SceneAsset)","fullName":"AdvancedSceneManager.Utility.SceneUtility.FindASMScene(UnityEditor.SceneAsset)","nameWithType":"SceneUtility.FindASMScene(SceneAsset)"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes*","name":"GetAllOpenUnityScenes","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_GetAllOpenUnityScenes_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.GetAllOpenUnityScenes","nameWithType":"SceneUtility.GetAllOpenUnityScenes"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.isStartupScene*","name":"isStartupScene","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_isStartupScene_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.isStartupScene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.isStartupScene","nameWithType":"SceneUtility.isStartupScene"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes*","name":"hasAnyScenes","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_hasAnyScenes_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.hasAnyScenes","nameWithType":"SceneUtility.hasAnyScenes"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.sceneCount*","name":"sceneCount","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_sceneCount_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.sceneCount","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.sceneCount","nameWithType":"SceneUtility.sceneCount"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Move*","name":"Move","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Move_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.Move","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.Move","nameWithType":"SceneUtility.Move"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.CreateDynamic*","name":"CreateDynamic","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_CreateDynamic_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.CreateDynamic","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.CreateDynamic","nameWithType":"SceneUtility.CreateDynamic"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder*","name":"CreateInCurrentFolder","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_CreateInCurrentFolder_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.CreateInCurrentFolder","nameWithType":"SceneUtility.CreateInCurrentFolder"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Create*","name":"Create","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Create_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.Create","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.Create","nameWithType":"SceneUtility.Create"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Remove_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.Remove","nameWithType":"SceneUtility.Remove"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.FindOpen*","name":"FindOpen","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_FindOpen_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.FindOpen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.FindOpen","nameWithType":"SceneUtility.FindOpen"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Find_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.Find","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.Find","nameWithType":"SceneUtility.Find"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene*","name":"MoveToNewScene","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_MoveToNewScene_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.MoveToNewScene","nameWithType":"SceneUtility.MoveToNewScene"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.MergeScenes*","name":"MergeScenes","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_MergeScenes_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.MergeScenes","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.MergeScenes","nameWithType":"SceneUtility.MergeScenes"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.Scene*","name":"Scene","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_Scene_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.Scene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.Scene","nameWithType":"SceneUtility.Scene"},{"uid":"AdvancedSceneManager.Utility.SceneUtility.FindASMScene*","name":"FindASMScene","href":"~/api/AdvancedSceneManager.Utility.SceneUtility.yml#AdvancedSceneManager_Utility_SceneUtility_FindASMScene_","commentId":"Overload:AdvancedSceneManager.Utility.SceneUtility.FindASMScene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SceneUtility.FindASMScene","nameWithType":"SceneUtility.FindASMScene"}],"api/AdvancedSceneManager.Callbacks.ICollectionClose.yml":[{"uid":"AdvancedSceneManager.Callbacks.ICollectionClose","name":"ICollectionClose","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionClose.yml","commentId":"T:AdvancedSceneManager.Callbacks.ICollectionClose","fullName":"AdvancedSceneManager.Callbacks.ICollectionClose","nameWithType":"ICollectionClose"},{"uid":"AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose(AdvancedSceneManager.Models.SceneCollection)","name":"OnCollectionClose(SceneCollection)","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionClose.yml#AdvancedSceneManager_Callbacks_ICollectionClose_OnCollectionClose_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ICollectionClose.OnCollectionClose(SceneCollection)"},{"uid":"AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose*","name":"OnCollectionClose","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionClose.yml#AdvancedSceneManager_Callbacks_ICollectionClose_OnCollectionClose_","commentId":"Overload:AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.ICollectionClose.OnCollectionClose","nameWithType":"ICollectionClose.OnCollectionClose"}],"api/AdvancedSceneManager.Callbacks.ParallelASMCallbacks.yml":[{"uid":"AdvancedSceneManager.Callbacks.ParallelASMCallbacks","name":"ParallelASMCallbacks","href":"~/api/AdvancedSceneManager.Callbacks.ParallelASMCallbacks.yml","commentId":"T:AdvancedSceneManager.Callbacks.ParallelASMCallbacks","fullName":"AdvancedSceneManager.Callbacks.ParallelASMCallbacks","nameWithType":"ParallelASMCallbacks"}],"api/AdvancedSceneManager.Core.Actions.AggregateAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction","name":"AggregateAction","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.AggregateAction","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction","nameWithType":"AggregateAction"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress","nameWithType":"AggregateAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.actions","name":"actions","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_actions","commentId":"P:AdvancedSceneManager.Core.Actions.AggregateAction.actions","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.actions","nameWithType":"AggregateAction.actions"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.#ctor(AdvancedSceneManager.Core.Actions.SceneAction[])","name":"AggregateAction(SceneAction[])","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction__ctor_AdvancedSceneManager_Core_Actions_SceneAction___","commentId":"M:AdvancedSceneManager.Core.Actions.AggregateAction.#ctor(AdvancedSceneManager.Core.Actions.SceneAction[])","name.vb":"AggregateAction(SceneAction())","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.AggregateAction(AdvancedSceneManager.Core.Actions.SceneAction[])","fullName.vb":"AdvancedSceneManager.Core.Actions.AggregateAction.AggregateAction(AdvancedSceneManager.Core.Actions.SceneAction())","nameWithType":"AggregateAction.AggregateAction(SceneAction[])","nameWithType.vb":"AggregateAction.AggregateAction(SceneAction())"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.#ctor(System.Action,AdvancedSceneManager.Core.Actions.SceneAction[])","name":"AggregateAction(Action, SceneAction[])","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction__ctor_System_Action_AdvancedSceneManager_Core_Actions_SceneAction___","commentId":"M:AdvancedSceneManager.Core.Actions.AggregateAction.#ctor(System.Action,AdvancedSceneManager.Core.Actions.SceneAction[])","name.vb":"AggregateAction(Action, SceneAction())","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.AggregateAction(System.Action, AdvancedSceneManager.Core.Actions.SceneAction[])","fullName.vb":"AdvancedSceneManager.Core.Actions.AggregateAction.AggregateAction(System.Action, AdvancedSceneManager.Core.Actions.SceneAction())","nameWithType":"AggregateAction.AggregateAction(Action, SceneAction[])","nameWithType.vb":"AggregateAction.AggregateAction(Action, SceneAction())"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.AggregateAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"AggregateAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.OnDone","name":"OnDone()","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_OnDone","commentId":"M:AdvancedSceneManager.Core.Actions.AggregateAction.OnDone","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.OnDone()","nameWithType":"AggregateAction.OnDone()"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.reportsProgress","nameWithType":"AggregateAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.actions*","name":"actions","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_actions_","commentId":"Overload:AdvancedSceneManager.Core.Actions.AggregateAction.actions","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.actions","nameWithType":"AggregateAction.actions"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.#ctor*","name":"AggregateAction","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.AggregateAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.AggregateAction","nameWithType":"AggregateAction.AggregateAction"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.AggregateAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.DoAction","nameWithType":"AggregateAction.DoAction"},{"uid":"AdvancedSceneManager.Core.Actions.AggregateAction.OnDone*","name":"OnDone","href":"~/api/AdvancedSceneManager.Core.Actions.AggregateAction.yml#AdvancedSceneManager_Core_Actions_AggregateAction_OnDone_","commentId":"Overload:AdvancedSceneManager.Core.Actions.AggregateAction.OnDone","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.AggregateAction.OnDone","nameWithType":"AggregateAction.OnDone"}],"api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction","name":"PlaySplashScreenAction","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction","nameWithType":"PlaySplashScreenAction"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress","nameWithType":"PlaySplashScreenAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.#ctor(System.Func{System.Collections.IEnumerator})","name":"PlaySplashScreenAction(Func<IEnumerator>)","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction__ctor_System_Func_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.#ctor(System.Func{System.Collections.IEnumerator})","name.vb":"PlaySplashScreenAction(Func(Of IEnumerator))","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.PlaySplashScreenAction(System.Func<System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.PlaySplashScreenAction(System.Func(Of System.Collections.IEnumerator))","nameWithType":"PlaySplashScreenAction.PlaySplashScreenAction(Func<IEnumerator>)","nameWithType.vb":"PlaySplashScreenAction.PlaySplashScreenAction(Func(Of IEnumerator))"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"PlaySplashScreenAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.reportsProgress","nameWithType":"PlaySplashScreenAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.#ctor*","name":"PlaySplashScreenAction","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.PlaySplashScreenAction","nameWithType":"PlaySplashScreenAction.PlaySplashScreenAction"},{"uid":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.yml#AdvancedSceneManager_Core_Actions_PlaySplashScreenAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.PlaySplashScreenAction.DoAction","nameWithType":"PlaySplashScreenAction.DoAction"}],"api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction","name":"SceneCloseCallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction","nameWithType":"SceneCloseCallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","name":"SceneCloseCallbackAction(OpenSceneInfo, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction__ctor_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.SceneCloseCallbackAction(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCloseCallbackAction.SceneCloseCallbackAction(OpenSceneInfo, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name":"SceneCloseCallbackAction(Func<OpenSceneInfo>, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction__ctor_System_Func_AdvancedSceneManager_Core_OpenSceneInfo__AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name.vb":"SceneCloseCallbackAction(Func(Of OpenSceneInfo), SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.SceneCloseCallbackAction(System.Func<AdvancedSceneManager.Core.OpenSceneInfo>, AdvancedSceneManager.Models.SceneCollection)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.SceneCloseCallbackAction(System.Func(Of AdvancedSceneManager.Core.OpenSceneInfo), AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCloseCallbackAction.SceneCloseCallbackAction(Func<OpenSceneInfo>, SceneCollection)","nameWithType.vb":"SceneCloseCallbackAction.SceneCloseCallbackAction(Func(Of OpenSceneInfo), SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction(ByRef System.Boolean)","nameWithType":"SceneCloseCallbackAction.BeforeDoAction(out Boolean)","nameWithType.vb":"SceneCloseCallbackAction.BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneCloseCallbackAction.DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor*","name":"SceneCloseCallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.SceneCloseCallbackAction","nameWithType":"SceneCloseCallbackAction.SceneCloseCallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.BeforeDoAction","nameWithType":"SceneCloseCallbackAction.BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseCallbackAction_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseCallbackAction.DoNonOverridenAction","nameWithType":"SceneCloseCallbackAction.DoNonOverridenAction"}],"api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction","name":"SceneOpenCallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction","nameWithType":"SceneOpenCallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","name":"SceneOpenCallbackAction(OpenSceneInfo, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction__ctor_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.SceneOpenCallbackAction(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneOpenCallbackAction.SceneOpenCallbackAction(OpenSceneInfo, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name":"SceneOpenCallbackAction(Func<OpenSceneInfo>, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction__ctor_System_Func_AdvancedSceneManager_Core_OpenSceneInfo__AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor(System.Func{AdvancedSceneManager.Core.OpenSceneInfo},AdvancedSceneManager.Models.SceneCollection)","name.vb":"SceneOpenCallbackAction(Func(Of OpenSceneInfo), SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.SceneOpenCallbackAction(System.Func<AdvancedSceneManager.Core.OpenSceneInfo>, AdvancedSceneManager.Models.SceneCollection)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.SceneOpenCallbackAction(System.Func(Of AdvancedSceneManager.Core.OpenSceneInfo), AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneOpenCallbackAction.SceneOpenCallbackAction(Func<OpenSceneInfo>, SceneCollection)","nameWithType.vb":"SceneOpenCallbackAction.SceneOpenCallbackAction(Func(Of OpenSceneInfo), SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction(ByRef System.Boolean)","nameWithType":"SceneOpenCallbackAction.BeforeDoAction(out Boolean)","nameWithType.vb":"SceneOpenCallbackAction.BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"SceneOpenCallbackAction.DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor*","name":"SceneOpenCallbackAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.SceneOpenCallbackAction","nameWithType":"SceneOpenCallbackAction.SceneOpenCallbackAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.BeforeDoAction","nameWithType":"SceneOpenCallbackAction.BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenCallbackAction_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenCallbackAction.DoNonOverridenAction","nameWithType":"SceneOpenCallbackAction.DoNonOverridenAction"}],"api/AdvancedSceneManager.Editor.Popup.yml":[{"uid":"AdvancedSceneManager.Editor.Popup","name":"Popup","href":"~/api/AdvancedSceneManager.Editor.Popup.yml","commentId":"T:AdvancedSceneManager.Editor.Popup","fullName":"AdvancedSceneManager.Editor.Popup","nameWithType":"Popup"},{"uid":"AdvancedSceneManager.Editor.Popup.OnClosed","name":"OnClosed","href":"~/api/AdvancedSceneManager.Editor.Popup.yml#AdvancedSceneManager_Editor_Popup_OnClosed","commentId":"E:AdvancedSceneManager.Editor.Popup.OnClosed","fullName":"AdvancedSceneManager.Editor.Popup.OnClosed","nameWithType":"Popup.OnClosed"},{"uid":"AdvancedSceneManager.Editor.Popup.RaiseOnClosed","name":"RaiseOnClosed()","href":"~/api/AdvancedSceneManager.Editor.Popup.yml#AdvancedSceneManager_Editor_Popup_RaiseOnClosed","commentId":"M:AdvancedSceneManager.Editor.Popup.RaiseOnClosed","fullName":"AdvancedSceneManager.Editor.Popup.RaiseOnClosed()","nameWithType":"Popup.RaiseOnClosed()"},{"uid":"AdvancedSceneManager.Editor.Popup.Reopen","name":"Reopen()","href":"~/api/AdvancedSceneManager.Editor.Popup.yml#AdvancedSceneManager_Editor_Popup_Reopen","commentId":"M:AdvancedSceneManager.Editor.Popup.Reopen","fullName":"AdvancedSceneManager.Editor.Popup.Reopen()","nameWithType":"Popup.Reopen()"},{"uid":"AdvancedSceneManager.Editor.Popup.RaiseOnClosed*","name":"RaiseOnClosed","href":"~/api/AdvancedSceneManager.Editor.Popup.yml#AdvancedSceneManager_Editor_Popup_RaiseOnClosed_","commentId":"Overload:AdvancedSceneManager.Editor.Popup.RaiseOnClosed","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup.RaiseOnClosed","nameWithType":"Popup.RaiseOnClosed"},{"uid":"AdvancedSceneManager.Editor.Popup.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Editor.Popup.yml#AdvancedSceneManager_Editor_Popup_Reopen_","commentId":"Overload:AdvancedSceneManager.Editor.Popup.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup.Reopen","nameWithType":"Popup.Reopen"}],"api/AdvancedSceneManager.Editor.SceneField.yml":[{"uid":"AdvancedSceneManager.Editor.SceneField","name":"SceneField","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml","commentId":"T:AdvancedSceneManager.Editor.SceneField","fullName":"AdvancedSceneManager.Editor.SceneField","nameWithType":"SceneField"},{"uid":"AdvancedSceneManager.Editor.SceneField.#ctor","name":"SceneField()","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField__ctor","commentId":"M:AdvancedSceneManager.Editor.SceneField.#ctor","fullName":"AdvancedSceneManager.Editor.SceneField.SceneField()","nameWithType":"SceneField.SceneField()"},{"uid":"AdvancedSceneManager.Editor.SceneField.labelFilter","name":"labelFilter","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_labelFilter","commentId":"P:AdvancedSceneManager.Editor.SceneField.labelFilter","fullName":"AdvancedSceneManager.Editor.SceneField.labelFilter","nameWithType":"SceneField.labelFilter"},{"uid":"AdvancedSceneManager.Editor.SceneField.showOpenButtons","name":"showOpenButtons","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_showOpenButtons","commentId":"P:AdvancedSceneManager.Editor.SceneField.showOpenButtons","fullName":"AdvancedSceneManager.Editor.SceneField.showOpenButtons","nameWithType":"SceneField.showOpenButtons"},{"uid":"AdvancedSceneManager.Editor.SceneField.defaultName","name":"defaultName","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_defaultName","commentId":"P:AdvancedSceneManager.Editor.SceneField.defaultName","fullName":"AdvancedSceneManager.Editor.SceneField.defaultName","nameWithType":"SceneField.defaultName"},{"uid":"AdvancedSceneManager.Editor.SceneField.Collection","name":"Collection","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_Collection","commentId":"P:AdvancedSceneManager.Editor.SceneField.Collection","fullName":"AdvancedSceneManager.Editor.SceneField.Collection","nameWithType":"SceneField.Collection"},{"uid":"AdvancedSceneManager.Editor.SceneField.OnSceneOpen","name":"OnSceneOpen","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_OnSceneOpen","commentId":"E:AdvancedSceneManager.Editor.SceneField.OnSceneOpen","fullName":"AdvancedSceneManager.Editor.SceneField.OnSceneOpen","nameWithType":"SceneField.OnSceneOpen"},{"uid":"AdvancedSceneManager.Editor.SceneField.OnSceneOpenAdditive","name":"OnSceneOpenAdditive","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_OnSceneOpenAdditive","commentId":"E:AdvancedSceneManager.Editor.SceneField.OnSceneOpenAdditive","fullName":"AdvancedSceneManager.Editor.SceneField.OnSceneOpenAdditive","nameWithType":"SceneField.OnSceneOpenAdditive"},{"uid":"AdvancedSceneManager.Editor.SceneField.OpenScene(AdvancedSceneManager.Models.Scene,System.Boolean,AdvancedSceneManager.Models.SceneCollection)","name":"OpenScene(Scene, Boolean, SceneCollection)","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_OpenScene_AdvancedSceneManager_Models_Scene_System_Boolean_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Editor.SceneField.OpenScene(AdvancedSceneManager.Models.Scene,System.Boolean,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Editor.SceneField.OpenScene(AdvancedSceneManager.Models.Scene, System.Boolean, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneField.OpenScene(Scene, Boolean, SceneCollection)"},{"uid":"AdvancedSceneManager.Editor.SceneField.onValueChanged","name":"onValueChanged","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_onValueChanged","commentId":"F:AdvancedSceneManager.Editor.SceneField.onValueChanged","fullName":"AdvancedSceneManager.Editor.SceneField.onValueChanged","nameWithType":"SceneField.onValueChanged"},{"uid":"AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify(AdvancedSceneManager.Models.Scene)","name":"SetValueWithoutNotify(Scene)","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_SetValueWithoutNotify_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify(AdvancedSceneManager.Models.Scene)","nameWithType":"SceneField.SetValueWithoutNotify(Scene)"},{"uid":"AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback(UnityEngine.UIElements.EventCallback{UnityEngine.UIElements.ChangeEvent{AdvancedSceneManager.Models.Scene}})","name":"RegisterValueChangedCallback(EventCallback<ChangeEvent<Scene>>)","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_RegisterValueChangedCallback_UnityEngine_UIElements_EventCallback_UnityEngine_UIElements_ChangeEvent_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback(UnityEngine.UIElements.EventCallback{UnityEngine.UIElements.ChangeEvent{AdvancedSceneManager.Models.Scene}})","name.vb":"RegisterValueChangedCallback(EventCallback(Of ChangeEvent(Of Scene)))","fullName":"AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback(UnityEngine.UIElements.EventCallback<UnityEngine.UIElements.ChangeEvent<AdvancedSceneManager.Models.Scene>>)","fullName.vb":"AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback(UnityEngine.UIElements.EventCallback(Of UnityEngine.UIElements.ChangeEvent(Of AdvancedSceneManager.Models.Scene)))","nameWithType":"SceneField.RegisterValueChangedCallback(EventCallback<ChangeEvent<Scene>>)","nameWithType.vb":"SceneField.RegisterValueChangedCallback(EventCallback(Of ChangeEvent(Of Scene)))"},{"uid":"AdvancedSceneManager.Editor.SceneField.value","name":"value","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_value","commentId":"P:AdvancedSceneManager.Editor.SceneField.value","fullName":"AdvancedSceneManager.Editor.SceneField.value","nameWithType":"SceneField.value"},{"uid":"AdvancedSceneManager.Editor.SceneField.#ctor*","name":"SceneField","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField__ctor_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.SceneField","nameWithType":"SceneField.SceneField"},{"uid":"AdvancedSceneManager.Editor.SceneField.labelFilter*","name":"labelFilter","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_labelFilter_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.labelFilter","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.labelFilter","nameWithType":"SceneField.labelFilter"},{"uid":"AdvancedSceneManager.Editor.SceneField.showOpenButtons*","name":"showOpenButtons","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_showOpenButtons_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.showOpenButtons","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.showOpenButtons","nameWithType":"SceneField.showOpenButtons"},{"uid":"AdvancedSceneManager.Editor.SceneField.defaultName*","name":"defaultName","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_defaultName_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.defaultName","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.defaultName","nameWithType":"SceneField.defaultName"},{"uid":"AdvancedSceneManager.Editor.SceneField.Collection*","name":"Collection","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_Collection_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.Collection","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.Collection","nameWithType":"SceneField.Collection"},{"uid":"AdvancedSceneManager.Editor.SceneField.OpenScene*","name":"OpenScene","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_OpenScene_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.OpenScene","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.OpenScene","nameWithType":"SceneField.OpenScene"},{"uid":"AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify*","name":"SetValueWithoutNotify","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_SetValueWithoutNotify_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.SetValueWithoutNotify","nameWithType":"SceneField.SetValueWithoutNotify"},{"uid":"AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback*","name":"RegisterValueChangedCallback","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_RegisterValueChangedCallback_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.RegisterValueChangedCallback","nameWithType":"SceneField.RegisterValueChangedCallback"},{"uid":"AdvancedSceneManager.Editor.SceneField.value*","name":"value","href":"~/api/AdvancedSceneManager.Editor.SceneField.yml#AdvancedSceneManager_Editor_SceneField_value_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.value","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.value","nameWithType":"SceneField.value"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement","name":"SceneManagerWindow.DragAndDropReorder.DragElement","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.list","name":"list","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_list","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.list","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.list","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.list"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.item","name":"item","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_item","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.item","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.item","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.item"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.button","name":"button","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_button","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.button","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.button","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.button"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseDown","name":"mouseDown","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_mouseDown","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseDown","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseDown","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.mouseDown"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseUp","name":"mouseUp","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_mouseUp","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseUp","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseUp","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.mouseUp"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseMove","name":"mouseMove","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_mouseMove","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseMove","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.mouseMove","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.mouseMove"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.index","name":"index","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_index","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.index","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.index","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.index"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootName","name":"itemRootName","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_itemRootName","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootName","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootName","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.itemRootName"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootClass","name":"itemRootClass","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_itemRootClass","commentId":"F:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootClass","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement.itemRootClass","nameWithType":"SceneManagerWindow.DragAndDropReorder.DragElement.itemRootClass"}],"api/AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility","name":"AssetsSavedUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.AssetsSavedUtility","fullName":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility","nameWithType":"AssetsSavedUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved","name":"onAssetsSaved","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.yml#AdvancedSceneManager_Editor_Utility_AssetsSavedUtility_onAssetsSaved","commentId":"E:AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved","fullName":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved","nameWithType":"AssetsSavedUtility.onAssetsSaved"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved2","name":"onAssetsSaved2","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.yml#AdvancedSceneManager_Editor_Utility_AssetsSavedUtility_onAssetsSaved2","commentId":"E:AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved2","fullName":"AdvancedSceneManager.Editor.Utility.AssetsSavedUtility.onAssetsSaved2","nameWithType":"AssetsSavedUtility.onAssetsSaved2"}],"api/AdvancedSceneManager.Editor.Utility.BlacklistUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.BlacklistUtility","name":"BlacklistUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.BlacklistUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.BlacklistUtility","fullName":"AdvancedSceneManager.Editor.Utility.BlacklistUtility","nameWithType":"BlacklistUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked(System.String)","name":"IsBlocked(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.BlacklistUtility.yml#AdvancedSceneManager_Editor_Utility_BlacklistUtility_IsBlocked_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked(System.String)","nameWithType":"BlacklistUtility.IsBlocked(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked*","name":"IsBlocked","href":"~/api/AdvancedSceneManager.Editor.Utility.BlacklistUtility.yml#AdvancedSceneManager_Editor_Utility_BlacklistUtility_IsBlocked_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.BlacklistUtility.IsBlocked","nameWithType":"BlacklistUtility.IsBlocked"}],"api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper","name":"MenuItemHelper","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.MenuItemHelper","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper","nameWithType":"MenuItemHelper"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem","name":"InvokeThisMenuItem()","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_InvokeThisMenuItem","commentId":"M:AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem()","nameWithType":"MenuItemHelper.InvokeThisMenuItem()"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Action)","name":"Setup(MethodBase, Action)","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Setup_System_Reflection_MethodBase_System_Action_","commentId":"M:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Action)","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase, System.Action)","nameWithType":"MenuItemHelper.Setup(MethodBase, Action)"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Func{System.Boolean},System.Action{System.Boolean})","name":"Setup(MethodBase, Func<Boolean>, Action<Boolean>)","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Setup_System_Reflection_MethodBase_System_Func_System_Boolean__System_Action_System_Boolean__","commentId":"M:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Func{System.Boolean},System.Action{System.Boolean})","name.vb":"Setup(MethodBase, Func(Of Boolean), Action(Of Boolean))","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase, System.Func<System.Boolean>, System.Action<System.Boolean>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase, System.Func(Of System.Boolean), System.Action(Of System.Boolean))","nameWithType":"MenuItemHelper.Setup(MethodBase, Func<Boolean>, Action<Boolean>)","nameWithType.vb":"MenuItemHelper.Setup(MethodBase, Func(Of Boolean), Action(Of Boolean))"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Reflection.PropertyInfo,System.Action{System.Boolean},System.Object)","name":"Setup(MethodBase, PropertyInfo, Action<Boolean>, Object)","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Setup_System_Reflection_MethodBase_System_Reflection_PropertyInfo_System_Action_System_Boolean__System_Object_","commentId":"M:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase,System.Reflection.PropertyInfo,System.Action{System.Boolean},System.Object)","name.vb":"Setup(MethodBase, PropertyInfo, Action(Of Boolean), Object)","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase, System.Reflection.PropertyInfo, System.Action<System.Boolean>, System.Object)","fullName.vb":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup(System.Reflection.MethodBase, System.Reflection.PropertyInfo, System.Action(Of System.Boolean), System.Object)","nameWithType":"MenuItemHelper.Setup(MethodBase, PropertyInfo, Action<Boolean>, Object)","nameWithType.vb":"MenuItemHelper.Setup(MethodBase, PropertyInfo, Action(Of Boolean), Object)"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh","name":"Refresh()","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Refresh","commentId":"M:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh()","nameWithType":"MenuItemHelper.Refresh()"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem*","name":"InvokeThisMenuItem","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_InvokeThisMenuItem_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.InvokeThisMenuItem","nameWithType":"MenuItemHelper.InvokeThisMenuItem"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup*","name":"Setup","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Setup_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Setup","nameWithType":"MenuItemHelper.Setup"},{"uid":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh*","name":"Refresh","href":"~/api/AdvancedSceneManager.Editor.Utility.MenuItemHelper.yml#AdvancedSceneManager_Editor_Utility_MenuItemHelper_Refresh_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.MenuItemHelper.Refresh","nameWithType":"MenuItemHelper.Refresh"}],"api/AdvancedSceneManager.Editor.Utility.OnGUIPrompt.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt","name":"OnGUIPrompt","href":"~/api/AdvancedSceneManager.Editor.Utility.OnGUIPrompt.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.OnGUIPrompt","fullName":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt","nameWithType":"OnGUIPrompt"},{"uid":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent,System.Action,System.Action,System.Action,System.Action,System.Action,System.Boolean,System.Boolean,System.String,UnityEngine.RectOffset,System.Nullable{UnityEngine.Vector2})","name":"Prompt(GUIContent, Action, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable<Vector2>)","href":"~/api/AdvancedSceneManager.Editor.Utility.OnGUIPrompt.yml#AdvancedSceneManager_Editor_Utility_OnGUIPrompt_Prompt_UnityEngine_GUIContent_System_Action_System_Action_System_Action_System_Action_System_Action_System_Boolean_System_Boolean_System_String_UnityEngine_RectOffset_System_Nullable_UnityEngine_Vector2__","commentId":"M:AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent,System.Action,System.Action,System.Action,System.Action,System.Action,System.Boolean,System.Boolean,System.String,UnityEngine.RectOffset,System.Nullable{UnityEngine.Vector2})","name.vb":"Prompt(GUIContent, Action, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable(Of Vector2))","fullName":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent, System.Action, System.Action, System.Action, System.Action, System.Action, System.Boolean, System.Boolean, System.String, UnityEngine.RectOffset, System.Nullable<UnityEngine.Vector2>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent, System.Action, System.Action, System.Action, System.Action, System.Action, System.Boolean, System.Boolean, System.String, UnityEngine.RectOffset, System.Nullable(Of UnityEngine.Vector2))","nameWithType":"OnGUIPrompt.Prompt(GUIContent, Action, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable<Vector2>)","nameWithType.vb":"OnGUIPrompt.Prompt(GUIContent, Action, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable(Of Vector2))"},{"uid":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent,System.Action,System.Action{System.Boolean}@,System.Action{System.Boolean}@,System.Action,System.Action,System.Action,System.Action,System.Boolean,System.Boolean,System.String,UnityEngine.RectOffset,System.Nullable{UnityEngine.Vector2})","name":"Prompt(GUIContent, Action, out Action<Boolean>, out Action<Boolean>, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable<Vector2>)","href":"~/api/AdvancedSceneManager.Editor.Utility.OnGUIPrompt.yml#AdvancedSceneManager_Editor_Utility_OnGUIPrompt_Prompt_UnityEngine_GUIContent_System_Action_System_Action_System_Boolean___System_Action_System_Boolean___System_Action_System_Action_System_Action_System_Action_System_Boolean_System_Boolean_System_String_UnityEngine_RectOffset_System_Nullable_UnityEngine_Vector2__","commentId":"M:AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent,System.Action,System.Action{System.Boolean}@,System.Action{System.Boolean}@,System.Action,System.Action,System.Action,System.Action,System.Boolean,System.Boolean,System.String,UnityEngine.RectOffset,System.Nullable{UnityEngine.Vector2})","name.vb":"Prompt(GUIContent, Action, ByRef Action(Of Boolean), ByRef Action(Of Boolean), Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable(Of Vector2))","fullName":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent, System.Action, out System.Action<System.Boolean>, out System.Action<System.Boolean>, System.Action, System.Action, System.Action, System.Action, System.Boolean, System.Boolean, System.String, UnityEngine.RectOffset, System.Nullable<UnityEngine.Vector2>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt(UnityEngine.GUIContent, System.Action, ByRef System.Action(Of System.Boolean), ByRef System.Action(Of System.Boolean), System.Action, System.Action, System.Action, System.Action, System.Boolean, System.Boolean, System.String, UnityEngine.RectOffset, System.Nullable(Of UnityEngine.Vector2))","nameWithType":"OnGUIPrompt.Prompt(GUIContent, Action, out Action<Boolean>, out Action<Boolean>, Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable<Vector2>)","nameWithType.vb":"OnGUIPrompt.Prompt(GUIContent, Action, ByRef Action(Of Boolean), ByRef Action(Of Boolean), Action, Action, Action, Action, Boolean, Boolean, String, RectOffset, Nullable(Of Vector2))"},{"uid":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt*","name":"Prompt","href":"~/api/AdvancedSceneManager.Editor.Utility.OnGUIPrompt.yml#AdvancedSceneManager_Editor_Utility_OnGUIPrompt_Prompt_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.OnGUIPrompt.Prompt","nameWithType":"OnGUIPrompt.Prompt"}],"api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions","name":"StyleExtensions","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.StyleExtensions","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions","nameWithType":"StyleExtensions"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name":"SetBorderWidth(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetBorderWidth_UnityEngine_UIElements_IStyle_System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__","commentId":"M:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name.vb":"SetBorderWidth(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth(UnityEngine.UIElements.IStyle, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth(UnityEngine.UIElements.IStyle, System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single))","nameWithType":"StyleExtensions.SetBorderWidth(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","nameWithType.vb":"StyleExtensions.SetBorderWidth(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor(UnityEngine.UIElements.IStyle,System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color})","name":"SetBorderColor(IStyle, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>)","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetBorderColor_UnityEngine_UIElements_IStyle_System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__System_Nullable_UnityEngine_Color__","commentId":"M:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor(UnityEngine.UIElements.IStyle,System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color},System.Nullable{UnityEngine.Color})","name.vb":"SetBorderColor(IStyle, Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color))","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor(UnityEngine.UIElements.IStyle, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>, System.Nullable<UnityEngine.Color>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor(UnityEngine.UIElements.IStyle, System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color), System.Nullable(Of UnityEngine.Color))","nameWithType":"StyleExtensions.SetBorderColor(IStyle, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>, Nullable<Color>)","nameWithType.vb":"StyleExtensions.SetBorderColor(IStyle, Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color), Nullable(Of Color))"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name":"SetMargin(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetMargin_UnityEngine_UIElements_IStyle_System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__","commentId":"M:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name.vb":"SetMargin(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin(UnityEngine.UIElements.IStyle, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin(UnityEngine.UIElements.IStyle, System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single))","nameWithType":"StyleExtensions.SetMargin(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","nameWithType.vb":"StyleExtensions.SetMargin(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name":"SetPadding(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetPadding_UnityEngine_UIElements_IStyle_System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__System_Nullable_System_Single__","commentId":"M:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding(UnityEngine.UIElements.IStyle,System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single},System.Nullable{System.Single})","name.vb":"SetPadding(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding(UnityEngine.UIElements.IStyle, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>, System.Nullable<System.Single>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding(UnityEngine.UIElements.IStyle, System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single), System.Nullable(Of System.Single))","nameWithType":"StyleExtensions.SetPadding(IStyle, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>, Nullable<Single>)","nameWithType.vb":"StyleExtensions.SetPadding(IStyle, Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single), Nullable(Of Single))"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth*","name":"SetBorderWidth","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetBorderWidth_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderWidth","nameWithType":"StyleExtensions.SetBorderWidth"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor*","name":"SetBorderColor","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetBorderColor_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetBorderColor","nameWithType":"StyleExtensions.SetBorderColor"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin*","name":"SetMargin","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetMargin_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetMargin","nameWithType":"StyleExtensions.SetMargin"},{"uid":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding*","name":"SetPadding","href":"~/api/AdvancedSceneManager.Editor.Utility.StyleExtensions.yml#AdvancedSceneManager_Editor_Utility_StyleExtensions_SetPadding_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.StyleExtensions.SetPadding","nameWithType":"StyleExtensions.SetPadding"}],"api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility","name":"TrimUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.TrimUtility","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility","nameWithType":"TrimUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel(UnityEngine.UIElements.TextElement,System.String,System.Func{System.Single},System.Boolean)","name":"TrimLabel(TextElement, String, Func<Single>, Boolean)","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml#AdvancedSceneManager_Editor_Utility_TrimUtility_TrimLabel_UnityEngine_UIElements_TextElement_System_String_System_Func_System_Single__System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel(UnityEngine.UIElements.TextElement,System.String,System.Func{System.Single},System.Boolean)","name.vb":"TrimLabel(TextElement, String, Func(Of Single), Boolean)","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel(UnityEngine.UIElements.TextElement, System.String, System.Func<System.Single>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel(UnityEngine.UIElements.TextElement, System.String, System.Func(Of System.Single), System.Boolean)","nameWithType":"TrimUtility.TrimLabel(TextElement, String, Func<Single>, Boolean)","nameWithType.vb":"TrimUtility.TrimLabel(TextElement, String, Func(Of Single), Boolean)"},{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.String,UnityEngine.UIElements.TextElement)","name":"GetLength(String, TextElement)","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml#AdvancedSceneManager_Editor_Utility_TrimUtility_GetLength_System_String_UnityEngine_UIElements_TextElement_","commentId":"M:AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.String,UnityEngine.UIElements.TextElement)","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.String, UnityEngine.UIElements.TextElement)","nameWithType":"TrimUtility.GetLength(String, TextElement)"},{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.Char,UnityEngine.UIElements.TextElement)","name":"GetLength(Char, TextElement)","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml#AdvancedSceneManager_Editor_Utility_TrimUtility_GetLength_System_Char_UnityEngine_UIElements_TextElement_","commentId":"M:AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.Char,UnityEngine.UIElements.TextElement)","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength(System.Char, UnityEngine.UIElements.TextElement)","nameWithType":"TrimUtility.GetLength(Char, TextElement)"},{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel*","name":"TrimLabel","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml#AdvancedSceneManager_Editor_Utility_TrimUtility_TrimLabel_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility.TrimLabel","nameWithType":"TrimUtility.TrimLabel"},{"uid":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength*","name":"GetLength","href":"~/api/AdvancedSceneManager.Editor.Utility.TrimUtility.yml#AdvancedSceneManager_Editor_Utility_TrimUtility_GetLength_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.TrimUtility.GetLength","nameWithType":"TrimUtility.GetLength"}],"api/AdvancedSceneManager.Models.CollectionStartupOption.yml":[{"uid":"AdvancedSceneManager.Models.CollectionStartupOption","name":"CollectionStartupOption","href":"~/api/AdvancedSceneManager.Models.CollectionStartupOption.yml","commentId":"T:AdvancedSceneManager.Models.CollectionStartupOption","fullName":"AdvancedSceneManager.Models.CollectionStartupOption","nameWithType":"CollectionStartupOption"},{"uid":"AdvancedSceneManager.Models.CollectionStartupOption.Auto","name":"Auto","href":"~/api/AdvancedSceneManager.Models.CollectionStartupOption.yml#AdvancedSceneManager_Models_CollectionStartupOption_Auto","commentId":"F:AdvancedSceneManager.Models.CollectionStartupOption.Auto","fullName":"AdvancedSceneManager.Models.CollectionStartupOption.Auto","nameWithType":"CollectionStartupOption.Auto"},{"uid":"AdvancedSceneManager.Models.CollectionStartupOption.Open","name":"Open","href":"~/api/AdvancedSceneManager.Models.CollectionStartupOption.yml#AdvancedSceneManager_Models_CollectionStartupOption_Open","commentId":"F:AdvancedSceneManager.Models.CollectionStartupOption.Open","fullName":"AdvancedSceneManager.Models.CollectionStartupOption.Open","nameWithType":"CollectionStartupOption.Open"},{"uid":"AdvancedSceneManager.Models.CollectionStartupOption.OpenAsPersistent","name":"OpenAsPersistent","href":"~/api/AdvancedSceneManager.Models.CollectionStartupOption.yml#AdvancedSceneManager_Models_CollectionStartupOption_OpenAsPersistent","commentId":"F:AdvancedSceneManager.Models.CollectionStartupOption.OpenAsPersistent","fullName":"AdvancedSceneManager.Models.CollectionStartupOption.OpenAsPersistent","nameWithType":"CollectionStartupOption.OpenAsPersistent"},{"uid":"AdvancedSceneManager.Models.CollectionStartupOption.DoNotOpen","name":"DoNotOpen","href":"~/api/AdvancedSceneManager.Models.CollectionStartupOption.yml#AdvancedSceneManager_Models_CollectionStartupOption_DoNotOpen","commentId":"F:AdvancedSceneManager.Models.CollectionStartupOption.DoNotOpen","fullName":"AdvancedSceneManager.Models.CollectionStartupOption.DoNotOpen","nameWithType":"CollectionStartupOption.DoNotOpen"}],"api/AdvancedSceneManager.Models.CollectionThreadPriority.yml":[{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority","name":"CollectionThreadPriority","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml","commentId":"T:AdvancedSceneManager.Models.CollectionThreadPriority","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority","nameWithType":"CollectionThreadPriority"},{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority.Auto","name":"Auto","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml#AdvancedSceneManager_Models_CollectionThreadPriority_Auto","commentId":"F:AdvancedSceneManager.Models.CollectionThreadPriority.Auto","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority.Auto","nameWithType":"CollectionThreadPriority.Auto"},{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority.Low","name":"Low","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml#AdvancedSceneManager_Models_CollectionThreadPriority_Low","commentId":"F:AdvancedSceneManager.Models.CollectionThreadPriority.Low","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority.Low","nameWithType":"CollectionThreadPriority.Low"},{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority.BelowNormal","name":"BelowNormal","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml#AdvancedSceneManager_Models_CollectionThreadPriority_BelowNormal","commentId":"F:AdvancedSceneManager.Models.CollectionThreadPriority.BelowNormal","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority.BelowNormal","nameWithType":"CollectionThreadPriority.BelowNormal"},{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority.Normal","name":"Normal","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml#AdvancedSceneManager_Models_CollectionThreadPriority_Normal","commentId":"F:AdvancedSceneManager.Models.CollectionThreadPriority.Normal","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority.Normal","nameWithType":"CollectionThreadPriority.Normal"},{"uid":"AdvancedSceneManager.Models.CollectionThreadPriority.High","name":"High","href":"~/api/AdvancedSceneManager.Models.CollectionThreadPriority.yml#AdvancedSceneManager_Models_CollectionThreadPriority_High","commentId":"F:AdvancedSceneManager.Models.CollectionThreadPriority.High","fullName":"AdvancedSceneManager.Models.CollectionThreadPriority.High","nameWithType":"CollectionThreadPriority.High"}],"api/AdvancedSceneManager.Models.yml":[{"uid":"AdvancedSceneManager.Models","name":"AdvancedSceneManager.Models","href":"~/api/AdvancedSceneManager.Models.yml","commentId":"N:AdvancedSceneManager.Models","fullName":"AdvancedSceneManager.Models","nameWithType":"AdvancedSceneManager.Models"}],"api/AdvancedSceneManager.SceneManager.yml":[{"uid":"AdvancedSceneManager.SceneManager","name":"SceneManager","href":"~/api/AdvancedSceneManager.SceneManager.yml","commentId":"T:AdvancedSceneManager.SceneManager","fullName":"AdvancedSceneManager.SceneManager","nameWithType":"SceneManager"},{"uid":"AdvancedSceneManager.SceneManager.assetManagement","name":"assetManagement","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_assetManagement","commentId":"P:AdvancedSceneManager.SceneManager.assetManagement","fullName":"AdvancedSceneManager.SceneManager.assetManagement","nameWithType":"SceneManager.assetManagement"},{"uid":"AdvancedSceneManager.SceneManager.collection","name":"collection","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_collection","commentId":"P:AdvancedSceneManager.SceneManager.collection","fullName":"AdvancedSceneManager.SceneManager.collection","nameWithType":"SceneManager.collection"},{"uid":"AdvancedSceneManager.SceneManager.standalone","name":"standalone","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_standalone","commentId":"P:AdvancedSceneManager.SceneManager.standalone","fullName":"AdvancedSceneManager.SceneManager.standalone","nameWithType":"SceneManager.standalone"},{"uid":"AdvancedSceneManager.SceneManager.utility","name":"utility","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_utility","commentId":"P:AdvancedSceneManager.SceneManager.utility","fullName":"AdvancedSceneManager.SceneManager.utility","nameWithType":"SceneManager.utility"},{"uid":"AdvancedSceneManager.SceneManager.runtime","name":"runtime","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_runtime","commentId":"P:AdvancedSceneManager.SceneManager.runtime","fullName":"AdvancedSceneManager.SceneManager.runtime","nameWithType":"SceneManager.runtime"},{"uid":"AdvancedSceneManager.SceneManager.settings","name":"settings","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_settings","commentId":"P:AdvancedSceneManager.SceneManager.settings","fullName":"AdvancedSceneManager.SceneManager.settings","nameWithType":"SceneManager.settings"},{"uid":"AdvancedSceneManager.SceneManager.profile","name":"profile","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_profile","commentId":"P:AdvancedSceneManager.SceneManager.profile","fullName":"AdvancedSceneManager.SceneManager.profile","nameWithType":"SceneManager.profile"},{"uid":"AdvancedSceneManager.SceneManager.editor","name":"editor","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_editor","commentId":"P:AdvancedSceneManager.SceneManager.editor","fullName":"AdvancedSceneManager.SceneManager.editor","nameWithType":"SceneManager.editor"},{"uid":"AdvancedSceneManager.SceneManager.assetManagement*","name":"assetManagement","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_assetManagement_","commentId":"Overload:AdvancedSceneManager.SceneManager.assetManagement","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.assetManagement","nameWithType":"SceneManager.assetManagement"},{"uid":"AdvancedSceneManager.SceneManager.collection*","name":"collection","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_collection_","commentId":"Overload:AdvancedSceneManager.SceneManager.collection","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.collection","nameWithType":"SceneManager.collection"},{"uid":"AdvancedSceneManager.SceneManager.standalone*","name":"standalone","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_standalone_","commentId":"Overload:AdvancedSceneManager.SceneManager.standalone","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.standalone","nameWithType":"SceneManager.standalone"},{"uid":"AdvancedSceneManager.SceneManager.utility*","name":"utility","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_utility_","commentId":"Overload:AdvancedSceneManager.SceneManager.utility","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.utility","nameWithType":"SceneManager.utility"},{"uid":"AdvancedSceneManager.SceneManager.runtime*","name":"runtime","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_runtime_","commentId":"Overload:AdvancedSceneManager.SceneManager.runtime","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.runtime","nameWithType":"SceneManager.runtime"},{"uid":"AdvancedSceneManager.SceneManager.settings*","name":"settings","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_settings_","commentId":"Overload:AdvancedSceneManager.SceneManager.settings","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.settings","nameWithType":"SceneManager.settings"},{"uid":"AdvancedSceneManager.SceneManager.profile*","name":"profile","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_profile_","commentId":"Overload:AdvancedSceneManager.SceneManager.profile","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.profile","nameWithType":"SceneManager.profile"},{"uid":"AdvancedSceneManager.SceneManager.editor*","name":"editor","href":"~/api/AdvancedSceneManager.SceneManager.yml#AdvancedSceneManager_SceneManager_editor_","commentId":"Overload:AdvancedSceneManager.SceneManager.editor","isSpec":"True","fullName":"AdvancedSceneManager.SceneManager.editor","nameWithType":"SceneManager.editor"}],"api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml":[{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility","name":"InGameToolbarUtility","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml","commentId":"T:AdvancedSceneManager.Utility.InGameToolbarUtility","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility","nameWithType":"InGameToolbarUtility"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled","name":"isEnabled","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_isEnabled","commentId":"P:AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled","nameWithType":"InGameToolbarUtility.isEnabled"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault","name":"expandedByDefault","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_expandedByDefault","commentId":"P:AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault","nameWithType":"InGameToolbarUtility.expandedByDefault"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor","name":"isEnabledInEditor","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_isEnabledInEditor","commentId":"P:AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor","nameWithType":"InGameToolbarUtility.isEnabledInEditor"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled*","name":"isEnabled","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_isEnabled_","commentId":"Overload:AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled","isSpec":"True","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabled","nameWithType":"InGameToolbarUtility.isEnabled"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault*","name":"expandedByDefault","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_expandedByDefault_","commentId":"Overload:AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault","isSpec":"True","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.expandedByDefault","nameWithType":"InGameToolbarUtility.expandedByDefault"},{"uid":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor*","name":"isEnabledInEditor","href":"~/api/AdvancedSceneManager.Utility.InGameToolbarUtility.yml#AdvancedSceneManager_Utility_InGameToolbarUtility_isEnabledInEditor_","commentId":"Overload:AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor","isSpec":"True","fullName":"AdvancedSceneManager.Utility.InGameToolbarUtility.isEnabledInEditor","nameWithType":"InGameToolbarUtility.isEnabledInEditor"}],"api/AdvancedSceneManager.Utility.IQueueable.yml":[{"uid":"AdvancedSceneManager.Utility.IQueueable","name":"IQueueable","href":"~/api/AdvancedSceneManager.Utility.IQueueable.yml","commentId":"T:AdvancedSceneManager.Utility.IQueueable","fullName":"AdvancedSceneManager.Utility.IQueueable","nameWithType":"IQueueable"},{"uid":"AdvancedSceneManager.Utility.IQueueable.OnTurn(System.Action)","name":"OnTurn(Action)","href":"~/api/AdvancedSceneManager.Utility.IQueueable.yml#AdvancedSceneManager_Utility_IQueueable_OnTurn_System_Action_","commentId":"M:AdvancedSceneManager.Utility.IQueueable.OnTurn(System.Action)","fullName":"AdvancedSceneManager.Utility.IQueueable.OnTurn(System.Action)","nameWithType":"IQueueable.OnTurn(Action)"},{"uid":"AdvancedSceneManager.Utility.IQueueable.OnCancel","name":"OnCancel()","href":"~/api/AdvancedSceneManager.Utility.IQueueable.yml#AdvancedSceneManager_Utility_IQueueable_OnCancel","commentId":"M:AdvancedSceneManager.Utility.IQueueable.OnCancel","fullName":"AdvancedSceneManager.Utility.IQueueable.OnCancel()","nameWithType":"IQueueable.OnCancel()"},{"uid":"AdvancedSceneManager.Utility.IQueueable.OnTurn*","name":"OnTurn","href":"~/api/AdvancedSceneManager.Utility.IQueueable.yml#AdvancedSceneManager_Utility_IQueueable_OnTurn_","commentId":"Overload:AdvancedSceneManager.Utility.IQueueable.OnTurn","isSpec":"True","fullName":"AdvancedSceneManager.Utility.IQueueable.OnTurn","nameWithType":"IQueueable.OnTurn"},{"uid":"AdvancedSceneManager.Utility.IQueueable.OnCancel*","name":"OnCancel","href":"~/api/AdvancedSceneManager.Utility.IQueueable.yml#AdvancedSceneManager_Utility_IQueueable_OnCancel_","commentId":"Overload:AdvancedSceneManager.Utility.IQueueable.OnCancel","isSpec":"True","fullName":"AdvancedSceneManager.Utility.IQueueable.OnCancel","nameWithType":"IQueueable.OnCancel"}],"api/AdvancedSceneManager.Utility.SerializableStringBoolDict.yml":[{"uid":"AdvancedSceneManager.Utility.SerializableStringBoolDict","name":"SerializableStringBoolDict","href":"~/api/AdvancedSceneManager.Utility.SerializableStringBoolDict.yml","commentId":"T:AdvancedSceneManager.Utility.SerializableStringBoolDict","fullName":"AdvancedSceneManager.Utility.SerializableStringBoolDict","nameWithType":"SerializableStringBoolDict"}],"api/AdvancedSceneManager.Utility.TimeSpanUtility.yml":[{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility","name":"TimeSpanUtility","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml","commentId":"T:AdvancedSceneManager.Utility.TimeSpanUtility","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility","nameWithType":"TimeSpanUtility"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.TimeSpan,System.String)","name":"ToDisplayString(TimeSpan, String)","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_ToDisplayString_System_TimeSpan_System_String_","commentId":"M:AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.TimeSpan,System.String)","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.TimeSpan, System.String)","nameWithType":"TimeSpanUtility.ToDisplayString(TimeSpan, String)"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.Single,System.String)","name":"ToDisplayString(Single, String)","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_ToDisplayString_System_Single_System_String_","commentId":"M:AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.Single,System.String)","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString(System.Single, System.String)","nameWithType":"TimeSpanUtility.ToDisplayString(Single, String)"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components(System.TimeSpan,System.String)","name":"ToDisplayString_Components(TimeSpan, String)","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_ToDisplayString_Components_System_TimeSpan_System_String_","commentId":"M:AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components(System.TimeSpan,System.String)","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components(System.TimeSpan, System.String)","nameWithType":"TimeSpanUtility.ToDisplayString_Components(TimeSpan, String)"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components(System.Single,System.String)","name":"FormatUnits_Components(Single, String)","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_FormatUnits_Components_System_Single_System_String_","commentId":"M:AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components(System.Single,System.String)","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components(System.Single, System.String)","nameWithType":"TimeSpanUtility.FormatUnits_Components(Single, String)"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString*","name":"ToDisplayString","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_ToDisplayString_","commentId":"Overload:AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString","isSpec":"True","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString","nameWithType":"TimeSpanUtility.ToDisplayString"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components*","name":"ToDisplayString_Components","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_ToDisplayString_Components_","commentId":"Overload:AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components","isSpec":"True","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.ToDisplayString_Components","nameWithType":"TimeSpanUtility.ToDisplayString_Components"},{"uid":"AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components*","name":"FormatUnits_Components","href":"~/api/AdvancedSceneManager.Utility.TimeSpanUtility.yml#AdvancedSceneManager_Utility_TimeSpanUtility_FormatUnits_Components_","commentId":"Overload:AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components","isSpec":"True","fullName":"AdvancedSceneManager.Utility.TimeSpanUtility.FormatUnits_Components","nameWithType":"TimeSpanUtility.FormatUnits_Components"}],"api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml":[{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1","name":"CallbackUtility.FluentInvokeAPI<T>","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml","commentId":"T:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1","name.vb":"CallbackUtility.FluentInvokeAPI(Of T)","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T)","nameWithType":"CallbackUtility.FluentInvokeAPI<T>","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T)"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.hasDefaultCallback","name":"hasDefaultCallback","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_hasDefaultCallback","commentId":"P:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.hasDefaultCallback","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.hasDefaultCallback","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).hasDefaultCallback","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.hasDefaultCallback","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).hasDefaultCallback"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithCallback(System.Func{`0,System.Collections.IEnumerator})","name":"WithCallback(Func<T, IEnumerator>)","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_WithCallback_System_Func__0_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithCallback(System.Func{`0,System.Collections.IEnumerator})","name.vb":"WithCallback(Func(Of T, IEnumerator))","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.WithCallback(System.Func<T, System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).WithCallback(System.Func(Of T, System.Collections.IEnumerator))","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.WithCallback(Func<T, IEnumerator>)","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).WithCallback(Func(Of T, IEnumerator))"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithParam(System.Object)","name":"WithParam(Object)","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_WithParam_System_Object_","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithParam(System.Object)","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.WithParam(System.Object)","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).WithParam(System.Object)","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.WithParam(Object)","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).WithParam(Object)"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Models.Scene[])","name":"On(Scene[])","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_On_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Models.Scene[])","name.vb":"On(Scene())","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.On(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).On(AdvancedSceneManager.Models.Scene())","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.On(Scene[])","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).On(Scene())"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Scene[])","name":"On(SceneCollection, Scene[])","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_On_AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Scene[])","name.vb":"On(SceneCollection, Scene())","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.On(AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).On(AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Scene())","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.On(SceneCollection, Scene[])","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).On(SceneCollection, Scene())"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.OnAllOpenScenes","name":"OnAllOpenScenes()","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_OnAllOpenScenes","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.OnAllOpenScenes","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.OnAllOpenScenes()","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).OnAllOpenScenes()","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.OnAllOpenScenes()","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).OnAllOpenScenes()"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"On(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_On_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"On(OpenSceneInfo())","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.On(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).On(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.On(OpenSceneInfo[])","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).On(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.hasDefaultCallback*","name":"hasDefaultCallback","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_hasDefaultCallback_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.hasDefaultCallback","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.hasDefaultCallback","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).hasDefaultCallback","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.hasDefaultCallback","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).hasDefaultCallback"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithCallback*","name":"WithCallback","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_WithCallback_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithCallback","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.WithCallback","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).WithCallback","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.WithCallback","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).WithCallback"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithParam*","name":"WithParam","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_WithParam_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.WithParam","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.WithParam","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).WithParam","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.WithParam","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).WithParam"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On*","name":"On","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_On_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.On","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.On","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).On","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.On","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).On"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.OnAllOpenScenes*","name":"OnAllOpenScenes","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI-1.yml#AdvancedSceneManager_Callbacks_CallbackUtility_FluentInvokeAPI_1_OnAllOpenScenes_","commentId":"Overload:AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI`1.OnAllOpenScenes","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI<T>.OnAllOpenScenes","fullName.vb":"AdvancedSceneManager.Callbacks.CallbackUtility.FluentInvokeAPI(Of T).OnAllOpenScenes","nameWithType":"CallbackUtility.FluentInvokeAPI<T>.OnAllOpenScenes","nameWithType.vb":"CallbackUtility.FluentInvokeAPI(Of T).OnAllOpenScenes"}],"api/AdvancedSceneManager.Callbacks.ICollectionOpen.yml":[{"uid":"AdvancedSceneManager.Callbacks.ICollectionOpen","name":"ICollectionOpen","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionOpen.yml","commentId":"T:AdvancedSceneManager.Callbacks.ICollectionOpen","fullName":"AdvancedSceneManager.Callbacks.ICollectionOpen","nameWithType":"ICollectionOpen"},{"uid":"AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen(AdvancedSceneManager.Models.SceneCollection)","name":"OnCollectionOpen(SceneCollection)","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionOpen.yml#AdvancedSceneManager_Callbacks_ICollectionOpen_OnCollectionOpen_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ICollectionOpen.OnCollectionOpen(SceneCollection)"},{"uid":"AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen*","name":"OnCollectionOpen","href":"~/api/AdvancedSceneManager.Callbacks.ICollectionOpen.yml#AdvancedSceneManager_Callbacks_ICollectionOpen_OnCollectionOpen_","commentId":"Overload:AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.ICollectionOpen.OnCollectionOpen","nameWithType":"ICollectionOpen.OnCollectionOpen"}],"api/AdvancedSceneManager.Editor.SceneAssetEditor.yml":[{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor","name":"SceneAssetEditor","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml","commentId":"T:AdvancedSceneManager.Editor.SceneAssetEditor","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor","nameWithType":"SceneAssetEditor"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_rootVisualElement","commentId":"P:AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement","nameWithType":"SceneAssetEditor.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.position","name":"position","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_position","commentId":"P:AdvancedSceneManager.Editor.SceneAssetEditor.position","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.position","nameWithType":"SceneAssetEditor.position"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI","name":"OnHeaderGUI()","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_OnHeaderGUI","commentId":"M:AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI()","nameWithType":"SceneAssetEditor.OnHeaderGUI()"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI","name":"CreateInspectorGUI()","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_CreateInspectorGUI","commentId":"M:AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI()","nameWithType":"SceneAssetEditor.CreateInspectorGUI()"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement*","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_rootVisualElement_","commentId":"Overload:AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.rootVisualElement","nameWithType":"SceneAssetEditor.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.position*","name":"position","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_position_","commentId":"Overload:AdvancedSceneManager.Editor.SceneAssetEditor.position","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.position","nameWithType":"SceneAssetEditor.position"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI*","name":"OnHeaderGUI","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_OnHeaderGUI_","commentId":"Overload:AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.OnHeaderGUI","nameWithType":"SceneAssetEditor.OnHeaderGUI"},{"uid":"AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI*","name":"CreateInspectorGUI","href":"~/api/AdvancedSceneManager.Editor.SceneAssetEditor.yml#AdvancedSceneManager_Editor_SceneAssetEditor_CreateInspectorGUI_","commentId":"Overload:AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneAssetEditor.CreateInspectorGUI","nameWithType":"SceneAssetEditor.CreateInspectorGUI"}],"api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml":[{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder","name":"SceneManagerWindow.DragAndDropReorder","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml","commentId":"T:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder","nameWithType":"SceneManagerWindow.DragAndDropReorder"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_rootVisualElement","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement","nameWithType":"SceneManagerWindow.DragAndDropReorder.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragStarted","name":"OnDragStarted","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_OnDragStarted","commentId":"E:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragStarted","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragStarted","nameWithType":"SceneManagerWindow.DragAndDropReorder.OnDragStarted"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragEnded","name":"OnDragEnded","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_OnDragEnded","commentId":"E:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragEnded","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragEnded","nameWithType":"SceneManagerWindow.DragAndDropReorder.OnDragEnded"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragCancel","name":"OnDragCancel","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_OnDragCancel","commentId":"E:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragCancel","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.OnDragCancel","nameWithType":"SceneManagerWindow.DragAndDropReorder.OnDragCancel"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement","name":"currentDragElement","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_currentDragElement","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement","nameWithType":"SceneManagerWindow.DragAndDropReorder.currentDragElement"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex","name":"newIndex","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_newIndex","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex","nameWithType":"SceneManagerWindow.DragAndDropReorder.newIndex"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset","name":"offset","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_offset","commentId":"P:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset","nameWithType":"SceneManagerWindow.DragAndDropReorder.offset"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList(UnityEngine.UIElements.VisualElement,System.String,System.String,System.String,System.String)","name":"RegisterList(VisualElement, String, String, String, String)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_RegisterList_UnityEngine_UIElements_VisualElement_System_String_System_String_System_String_System_String_","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList(UnityEngine.UIElements.VisualElement,System.String,System.String,System.String,System.String)","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList(UnityEngine.UIElements.VisualElement, System.String, System.String, System.String, System.String)","nameWithType":"SceneManagerWindow.DragAndDropReorder.RegisterList(VisualElement, String, String, String, String)"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList(UnityEngine.UIElements.VisualElement)","name":"UnregisterList(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_UnregisterList_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList(UnityEngine.UIElements.VisualElement)","nameWithType":"SceneManagerWindow.DragAndDropReorder.UnregisterList(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll","name":"UnregisterListAll()","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_UnregisterListAll","commentId":"M:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll()","nameWithType":"SceneManagerWindow.DragAndDropReorder.UnregisterListAll()"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement*","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_rootVisualElement_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.rootVisualElement","nameWithType":"SceneManagerWindow.DragAndDropReorder.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement*","name":"currentDragElement","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_currentDragElement_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.currentDragElement","nameWithType":"SceneManagerWindow.DragAndDropReorder.currentDragElement"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex*","name":"newIndex","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_newIndex_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.newIndex","nameWithType":"SceneManagerWindow.DragAndDropReorder.newIndex"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset*","name":"offset","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_offset_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.offset","nameWithType":"SceneManagerWindow.DragAndDropReorder.offset"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList*","name":"RegisterList","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_RegisterList_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.RegisterList","nameWithType":"SceneManagerWindow.DragAndDropReorder.RegisterList"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList*","name":"UnregisterList","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_UnregisterList_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterList","nameWithType":"SceneManagerWindow.DragAndDropReorder.UnregisterList"},{"uid":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll*","name":"UnregisterListAll","href":"~/api/AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.yml#AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_UnregisterListAll_","commentId":"Overload:AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.UnregisterListAll","nameWithType":"SceneManagerWindow.DragAndDropReorder.UnregisterListAll"}],"api/AdvancedSceneManager.Editor.SettingsTab.yml":[{"uid":"AdvancedSceneManager.Editor.SettingsTab","name":"SettingsTab","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml","commentId":"T:AdvancedSceneManager.Editor.SettingsTab","fullName":"AdvancedSceneManager.Editor.SettingsTab","nameWithType":"SettingsTab"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.Settings","name":"Settings","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_Settings","commentId":"P:AdvancedSceneManager.Editor.SettingsTab.Settings","fullName":"AdvancedSceneManager.Editor.SettingsTab.Settings","nameWithType":"SettingsTab.Settings"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.OnEnable(UnityEngine.UIElements.VisualElement)","name":"OnEnable(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_OnEnable_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.SettingsTab.OnEnable(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.SettingsTab.OnEnable(UnityEngine.UIElements.VisualElement)","nameWithType":"SettingsTab.OnEnable(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.InitializeProfile(UnityEngine.UIElements.VisualElement,System.Action)","name":"InitializeProfile(VisualElement, Action)","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_InitializeProfile_UnityEngine_UIElements_VisualElement_System_Action_","commentId":"M:AdvancedSceneManager.Editor.SettingsTab.InitializeProfile(UnityEngine.UIElements.VisualElement,System.Action)","fullName":"AdvancedSceneManager.Editor.SettingsTab.InitializeProfile(UnityEngine.UIElements.VisualElement, System.Action)","nameWithType":"SettingsTab.InitializeProfile(VisualElement, Action)"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.Settings*","name":"Settings","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_Settings_","commentId":"Overload:AdvancedSceneManager.Editor.SettingsTab.Settings","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SettingsTab.Settings","nameWithType":"SettingsTab.Settings"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.SettingsTab.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SettingsTab.OnEnable","nameWithType":"SettingsTab.OnEnable"},{"uid":"AdvancedSceneManager.Editor.SettingsTab.InitializeProfile*","name":"InitializeProfile","href":"~/api/AdvancedSceneManager.Editor.SettingsTab.yml#AdvancedSceneManager_Editor_SettingsTab_InitializeProfile_","commentId":"Overload:AdvancedSceneManager.Editor.SettingsTab.InitializeProfile","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SettingsTab.InitializeProfile","nameWithType":"SettingsTab.InitializeProfile"}],"api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.BuildError.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.BuildError","name":"BuildEventsUtility.BuildError","href":"~/api/AdvancedSceneManager.Editor.Utility.BuildEventsUtility.BuildError.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.BuildEventsUtility.BuildError","fullName":"AdvancedSceneManager.Editor.Utility.BuildEventsUtility.BuildError","nameWithType":"BuildEventsUtility.BuildError"}],"api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt","name":"GenericPrompt","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.GenericPrompt","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt","nameWithType":"GenericPrompt"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt(System.String,System.String,System.String,System.String,System.Single)","name":"Prompt(String, String, String, String, Single)","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_Prompt_System_String_System_String_System_String_System_String_System_Single_","commentId":"M:AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt(System.String,System.String,System.String,System.String,System.Single)","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt(System.String, System.String, System.String, System.String, System.Single)","nameWithType":"GenericPrompt.Prompt(String, String, String, String, Single)"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_extraHeight","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight","nameWithType":"GenericPrompt.extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.width","name":"width","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_width","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt.width","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.width","nameWithType":"GenericPrompt.width"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_title","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt.title","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.title","nameWithType":"GenericPrompt.title"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton","name":"cancelButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_cancelButton","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton","nameWithType":"GenericPrompt.cancelButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton","name":"okButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_okButton","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton","nameWithType":"GenericPrompt.okButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI(System.Object@)","name":"OnContentGUI(ref Object)","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_OnContentGUI_System_Object__","commentId":"M:AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI(System.Object@)","name.vb":"OnContentGUI(ByRef Object)","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI(ref System.Object)","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI(ByRef System.Object)","nameWithType":"GenericPrompt.OnContentGUI(ref Object)","nameWithType.vb":"GenericPrompt.OnContentGUI(ByRef Object)"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt*","name":"Prompt","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_Prompt_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.Prompt","nameWithType":"GenericPrompt.Prompt"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight*","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_extraHeight_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.extraHeight","nameWithType":"GenericPrompt.extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.width*","name":"width","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_width_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.width","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.width","nameWithType":"GenericPrompt.width"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.title","nameWithType":"GenericPrompt.title"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton*","name":"cancelButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_cancelButton_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.cancelButton","nameWithType":"GenericPrompt.cancelButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton*","name":"okButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_okButton_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.okButton","nameWithType":"GenericPrompt.okButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt.OnContentGUI","nameWithType":"GenericPrompt.OnContentGUI"}],"api/AdvancedSceneManager.Editor.Utility.ListUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility","name":"ListUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.ListUtility","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility","nameWithType":"ListUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp``1(``0[]@,``0)","name":"MoveUp<T>(ref T[], T)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_MoveUp__1___0______0_","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp``1(``0[]@,``0)","name.vb":"MoveUp(Of T)(ByRef T(), T)","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp<T>(ref T[], T)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp(Of T)(ByRef T(), T)","nameWithType":"ListUtility.MoveUp<T>(ref T[], T)","nameWithType.vb":"ListUtility.MoveUp(Of T)(ByRef T(), T)"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown``1(``0[]@,``0)","name":"MoveDown<T>(ref T[], T)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_MoveDown__1___0______0_","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown``1(``0[]@,``0)","name.vb":"MoveDown(Of T)(ByRef T(), T)","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown<T>(ref T[], T)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown(Of T)(ByRef T(), T)","nameWithType":"ListUtility.MoveDown<T>(ref T[], T)","nameWithType.vb":"ListUtility.MoveDown(Of T)(ByRef T(), T)"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach``1(``0[],System.Action{``0,System.Int32})","name":"ForEach<T>(T[], Action<T, Int32>)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_ForEach__1___0___System_Action___0_System_Int32__","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.ForEach``1(``0[],System.Action{``0,System.Int32})","name.vb":"ForEach(Of T)(T(), Action(Of T, Int32))","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach<T>(T[], System.Action<T, System.Int32>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach(Of T)(T(), System.Action(Of T, System.Int32))","nameWithType":"ListUtility.ForEach<T>(T[], Action<T, Int32>)","nameWithType.vb":"ListUtility.ForEach(Of T)(T(), Action(Of T, Int32))"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach``1(System.Collections.Generic.IEnumerable{``0},System.Action{``0,System.Int32})","name":"ForEach<T>(IEnumerable<T>, Action<T, Int32>)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_ForEach__1_System_Collections_Generic_IEnumerable___0__System_Action___0_System_Int32__","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.ForEach``1(System.Collections.Generic.IEnumerable{``0},System.Action{``0,System.Int32})","name.vb":"ForEach(Of T)(IEnumerable(Of T), Action(Of T, Int32))","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach<T>(System.Collections.Generic.IEnumerable<T>, System.Action<T, System.Int32>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach(Of T)(System.Collections.Generic.IEnumerable(Of T), System.Action(Of T, System.Int32))","nameWithType":"ListUtility.ForEach<T>(IEnumerable<T>, Action<T, Int32>)","nameWithType.vb":"ListUtility.ForEach(Of T)(IEnumerable(Of T), Action(Of T, Int32))"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.Flatten``1(System.Collections.Generic.IEnumerable{``0},System.Func{``0,System.Collections.Generic.IEnumerable{``0}})","name":"Flatten<T>(IEnumerable<T>, Func<T, IEnumerable<T>>)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_Flatten__1_System_Collections_Generic_IEnumerable___0__System_Func___0_System_Collections_Generic_IEnumerable___0___","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.Flatten``1(System.Collections.Generic.IEnumerable{``0},System.Func{``0,System.Collections.Generic.IEnumerable{``0}})","name.vb":"Flatten(Of T)(IEnumerable(Of T), Func(Of T, IEnumerable(Of T)))","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.Flatten<T>(System.Collections.Generic.IEnumerable<T>, System.Func<T, System.Collections.Generic.IEnumerable<T>>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.Flatten(Of T)(System.Collections.Generic.IEnumerable(Of T), System.Func(Of T, System.Collections.Generic.IEnumerable(Of T)))","nameWithType":"ListUtility.Flatten<T>(IEnumerable<T>, Func<T, IEnumerable<T>>)","nameWithType.vb":"ListUtility.Flatten(Of T)(IEnumerable(Of T), Func(Of T, IEnumerable(Of T)))"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.Except``1(System.Collections.Generic.IEnumerable{``0},``0)","name":"Except<T>(IEnumerable<T>, T)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_Except__1_System_Collections_Generic_IEnumerable___0____0_","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.Except``1(System.Collections.Generic.IEnumerable{``0},``0)","name.vb":"Except(Of T)(IEnumerable(Of T), T)","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.Except<T>(System.Collections.Generic.IEnumerable<T>, T)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.Except(Of T)(System.Collections.Generic.IEnumerable(Of T), T)","nameWithType":"ListUtility.Except<T>(IEnumerable<T>, T)","nameWithType.vb":"ListUtility.Except(Of T)(IEnumerable(Of T), T)"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive``1(System.Collections.Generic.IEnumerable{``0},System.Func{``0,``0,System.Boolean})","name":"GroupConsecutive<T>(IEnumerable<T>, Func<T, T, Boolean>)","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_GroupConsecutive__1_System_Collections_Generic_IEnumerable___0__System_Func___0___0_System_Boolean__","commentId":"M:AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive``1(System.Collections.Generic.IEnumerable{``0},System.Func{``0,``0,System.Boolean})","name.vb":"GroupConsecutive(Of T)(IEnumerable(Of T), Func(Of T, T, Boolean))","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive<T>(System.Collections.Generic.IEnumerable<T>, System.Func<T, T, System.Boolean>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive(Of T)(System.Collections.Generic.IEnumerable(Of T), System.Func(Of T, T, System.Boolean))","nameWithType":"ListUtility.GroupConsecutive<T>(IEnumerable<T>, Func<T, T, Boolean>)","nameWithType.vb":"ListUtility.GroupConsecutive(Of T)(IEnumerable(Of T), Func(Of T, T, Boolean))"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp*","name":"MoveUp","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_MoveUp_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveUp","nameWithType":"ListUtility.MoveUp"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown*","name":"MoveDown","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_MoveDown_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.MoveDown","nameWithType":"ListUtility.MoveDown"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach*","name":"ForEach","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_ForEach_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.ForEach","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.ForEach","nameWithType":"ListUtility.ForEach"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.Flatten*","name":"Flatten","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_Flatten_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.Flatten","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.Flatten","nameWithType":"ListUtility.Flatten"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.Except*","name":"Except","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_Except_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.Except","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.Except","nameWithType":"ListUtility.Except"},{"uid":"AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive*","name":"GroupConsecutive","href":"~/api/AdvancedSceneManager.Editor.Utility.ListUtility.yml#AdvancedSceneManager_Editor_Utility_ListUtility_GroupConsecutive_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.ListUtility.GroupConsecutive","nameWithType":"ListUtility.GroupConsecutive"}],"api/AdvancedSceneManager.Editor.Utility.PromptName.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PromptName","name":"PromptName","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptName.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PromptName","fullName":"AdvancedSceneManager.Editor.Utility.PromptName","nameWithType":"PromptName"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptName.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptName.yml#AdvancedSceneManager_Editor_Utility_PromptName_title","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptName.title","fullName":"AdvancedSceneManager.Editor.Utility.PromptName.title","nameWithType":"PromptName.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI(System.String@)","name":"OnContentGUI(ref String)","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptName.yml#AdvancedSceneManager_Editor_Utility_PromptName_OnContentGUI_System_String__","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI(System.String@)","name.vb":"OnContentGUI(ByRef String)","fullName":"AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI(ref System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI(ByRef System.String)","nameWithType":"PromptName.OnContentGUI(ref String)","nameWithType.vb":"PromptName.OnContentGUI(ByRef String)"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptName.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptName.yml#AdvancedSceneManager_Editor_Utility_PromptName_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptName.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptName.title","nameWithType":"PromptName.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptName.yml#AdvancedSceneManager_Editor_Utility_PromptName_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptName.OnContentGUI","nameWithType":"PromptName.OnContentGUI"}],"api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage","name":"PromptNameAndMessage","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage","nameWithType":"PromptNameAndMessage"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_title","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title","nameWithType":"PromptNameAndMessage.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_extraHeight","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight","nameWithType":"PromptNameAndMessage.extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI(System.ValueTuple{System.String,System.String}@)","name":"OnContentGUI(ref (String name, String message))","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_OnContentGUI_System_ValueTuple_System_String_System_String___","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI(System.ValueTuple{System.String,System.String}@)","name.vb":"OnContentGUI(ByRef (name As String, message As String)(Of String, String))","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI(ref System.ValueTuple<System.String, System.String>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI(ByRef System.ValueTuple(Of System.String, System.String))","nameWithType":"PromptNameAndMessage.OnContentGUI(ref (String name, String message))","nameWithType.vb":"PromptNameAndMessage.OnContentGUI(ByRef (name As String, message As String)(Of String, String))"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.title","nameWithType":"PromptNameAndMessage.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight*","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_extraHeight_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.extraHeight","nameWithType":"PromptNameAndMessage.extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.yml#AdvancedSceneManager_Editor_Utility_PromptNameAndMessage_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptNameAndMessage.OnContentGUI","nameWithType":"PromptNameAndMessage.OnContentGUI"}],"api/AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.yml":[{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction","name":"ASMSettings.Local.SaveAction","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.yml","commentId":"T:AdvancedSceneManager.Models.ASMSettings.Local.SaveAction","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction","nameWithType":"ASMSettings.Local.SaveAction"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.DoNothing","name":"DoNothing","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.yml#AdvancedSceneManager_Models_ASMSettings_Local_SaveAction_DoNothing","commentId":"F:AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.DoNothing","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.DoNothing","nameWithType":"ASMSettings.Local.SaveAction.DoNothing"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Save","name":"Save","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.yml#AdvancedSceneManager_Models_ASMSettings_Local_SaveAction_Save","commentId":"F:AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Save","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Save","nameWithType":"ASMSettings.Local.SaveAction.Save"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Prompt","name":"Prompt","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.yml#AdvancedSceneManager_Models_ASMSettings_Local_SaveAction_Prompt","commentId":"F:AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Prompt","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.SaveAction.Prompt","nameWithType":"ASMSettings.Local.SaveAction.Prompt"}],"api/AdvancedSceneManager.Models.ASMSettings.Local.yml":[{"uid":"AdvancedSceneManager.Models.ASMSettings.Local","name":"ASMSettings.Local","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml","commentId":"T:AdvancedSceneManager.Models.ASMSettings.Local","fullName":"AdvancedSceneManager.Models.ASMSettings.Local","nameWithType":"ASMSettings.Local"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild","name":"allowExcludingCollectionsFromBuild","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_allowExcludingCollectionsFromBuild","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild","nameWithType":"ASMSettings.Local.allowExcludingCollectionsFromBuild"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton","name":"displayCollectionPlayButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionPlayButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton","nameWithType":"ASMSettings.Local.displayCollectionPlayButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton","name":"displayCollectionOpenButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionOpenButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton","nameWithType":"ASMSettings.Local.displayCollectionOpenButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton","name":"displayCollectionAdditiveButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionAdditiveButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton","nameWithType":"ASMSettings.Local.displayCollectionAdditiveButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton","name":"displayExtraAddCollectionButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayExtraAddCollectionButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton","nameWithType":"ASMSettings.Local.displayExtraAddCollectionButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton","name":"displaySceneHelperDragButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displaySceneHelperDragButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton","nameWithType":"ASMSettings.Local.displaySceneHelperDragButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy","name":"displayPersistentIndicatorInHierarchy","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayPersistentIndicatorInHierarchy","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy","nameWithType":"ASMSettings.Local.displayPersistentIndicatorInHierarchy"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy","name":"displayCollectionTitleOnScenesInHierarchy","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionTitleOnScenesInHierarchy","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy","nameWithType":"ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections","name":"displayDynamicCollections","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayDynamicCollections","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections","nameWithType":"ASMSettings.Local.displayDynamicCollections"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings","name":"allowEditingOfBuildSettings","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_allowEditingOfBuildSettings","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings","nameWithType":"ASMSettings.Local.allowEditingOfBuildSettings"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated","name":"autoOpenScenesWhenCreated","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_autoOpenScenesWhenCreated","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated","nameWithType":"ASMSettings.Local.autoOpenScenesWhenCreated"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField","name":"useSaveDialogWhenCreatingScenesFromSceneField","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_useSaveDialogWhenCreatingScenesFromSceneField","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField","nameWithType":"ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen","name":"openAssociatedCollectionOnSceneAssetOpen","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_openAssociatedCollectionOnSceneAssetOpen","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen","nameWithType":"ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton","name":"saveActionWhenUsingASMPlayButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_saveActionWhenUsingASMPlayButton","commentId":"P:AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton","nameWithType":"ASMSettings.Local.saveActionWhenUsingASMPlayButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.Get``1(``0,System.String)","name":"Get<T>(T, String)","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_Get__1___0_System_String_","commentId":"M:AdvancedSceneManager.Models.ASMSettings.Local.Get``1(``0,System.String)","name.vb":"Get(Of T)(T, String)","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.Get<T>(T, System.String)","fullName.vb":"AdvancedSceneManager.Models.ASMSettings.Local.Get(Of T)(T, System.String)","nameWithType":"ASMSettings.Local.Get<T>(T, String)","nameWithType.vb":"ASMSettings.Local.Get(Of T)(T, String)"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.Set``1(``0,System.String)","name":"Set<T>(T, String)","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_Set__1___0_System_String_","commentId":"M:AdvancedSceneManager.Models.ASMSettings.Local.Set``1(``0,System.String)","name.vb":"Set(Of T)(T, String)","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.Set<T>(T, System.String)","fullName.vb":"AdvancedSceneManager.Models.ASMSettings.Local.Set(Of T)(T, System.String)","nameWithType":"ASMSettings.Local.Set<T>(T, String)","nameWithType.vb":"ASMSettings.Local.Set(Of T)(T, String)"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild*","name":"allowExcludingCollectionsFromBuild","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_allowExcludingCollectionsFromBuild_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.allowExcludingCollectionsFromBuild","nameWithType":"ASMSettings.Local.allowExcludingCollectionsFromBuild"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton*","name":"displayCollectionPlayButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionPlayButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionPlayButton","nameWithType":"ASMSettings.Local.displayCollectionPlayButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton*","name":"displayCollectionOpenButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionOpenButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionOpenButton","nameWithType":"ASMSettings.Local.displayCollectionOpenButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton*","name":"displayCollectionAdditiveButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionAdditiveButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionAdditiveButton","nameWithType":"ASMSettings.Local.displayCollectionAdditiveButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton*","name":"displayExtraAddCollectionButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayExtraAddCollectionButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayExtraAddCollectionButton","nameWithType":"ASMSettings.Local.displayExtraAddCollectionButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton*","name":"displaySceneHelperDragButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displaySceneHelperDragButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displaySceneHelperDragButton","nameWithType":"ASMSettings.Local.displaySceneHelperDragButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy*","name":"displayPersistentIndicatorInHierarchy","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayPersistentIndicatorInHierarchy_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayPersistentIndicatorInHierarchy","nameWithType":"ASMSettings.Local.displayPersistentIndicatorInHierarchy"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy*","name":"displayCollectionTitleOnScenesInHierarchy","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayCollectionTitleOnScenesInHierarchy_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy","nameWithType":"ASMSettings.Local.displayCollectionTitleOnScenesInHierarchy"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections*","name":"displayDynamicCollections","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_displayDynamicCollections_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.displayDynamicCollections","nameWithType":"ASMSettings.Local.displayDynamicCollections"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings*","name":"allowEditingOfBuildSettings","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_allowEditingOfBuildSettings_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.allowEditingOfBuildSettings","nameWithType":"ASMSettings.Local.allowEditingOfBuildSettings"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated*","name":"autoOpenScenesWhenCreated","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_autoOpenScenesWhenCreated_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.autoOpenScenesWhenCreated","nameWithType":"ASMSettings.Local.autoOpenScenesWhenCreated"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField*","name":"useSaveDialogWhenCreatingScenesFromSceneField","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_useSaveDialogWhenCreatingScenesFromSceneField_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField","nameWithType":"ASMSettings.Local.useSaveDialogWhenCreatingScenesFromSceneField"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen*","name":"openAssociatedCollectionOnSceneAssetOpen","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_openAssociatedCollectionOnSceneAssetOpen_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen","nameWithType":"ASMSettings.Local.openAssociatedCollectionOnSceneAssetOpen"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton*","name":"saveActionWhenUsingASMPlayButton","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_saveActionWhenUsingASMPlayButton_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.saveActionWhenUsingASMPlayButton","nameWithType":"ASMSettings.Local.saveActionWhenUsingASMPlayButton"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.Get*","name":"Get","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_Get_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.Get","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.Get","nameWithType":"ASMSettings.Local.Get"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Local.Set*","name":"Set","href":"~/api/AdvancedSceneManager.Models.ASMSettings.Local.yml#AdvancedSceneManager_Models_ASMSettings_Local_Set_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Local.Set","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Local.Set","nameWithType":"ASMSettings.Local.Set"}],"api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml":[{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate","name":"SceneCollectionTemplate","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml","commentId":"T:AdvancedSceneManager.Models.SceneCollectionTemplate","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate","nameWithType":"SceneCollectionTemplate"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.name","name":"name","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_name","commentId":"P:AdvancedSceneManager.Models.SceneCollectionTemplate.name","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.name","nameWithType":"SceneCollectionTemplate.name"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.title","name":"title","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_title","commentId":"P:AdvancedSceneManager.Models.SceneCollectionTemplate.title","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.title","nameWithType":"SceneCollectionTemplate.title"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection(AdvancedSceneManager.Models.Profile)","name":"CreateCollection(Profile)","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection(AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection(AdvancedSceneManager.Models.Profile)","nameWithType":"SceneCollectionTemplate.CreateCollection(Profile)"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.Apply(AdvancedSceneManager.Models.SceneCollection)","name":"Apply(SceneCollection)","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_Apply_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.SceneCollectionTemplate.Apply(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.Apply(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCollectionTemplate.Apply(SceneCollection)"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder(AdvancedSceneManager.Models.SceneCollection)","name":"CreateTemplateInCurrentFolder(SceneCollection)","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateTemplateInCurrentFolder_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCollectionTemplate.CreateTemplateInCurrentFolder(SceneCollection)"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate(System.String,AdvancedSceneManager.Models.SceneCollection)","name":"CreateTemplate(String, SceneCollection)","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateTemplate_System_String_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate(System.String,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate(System.String, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCollectionTemplate.CreateTemplate(String, SceneCollection)"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.name*","name":"name","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_name_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.name","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.name","nameWithType":"SceneCollectionTemplate.name"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.title*","name":"title","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_title_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.title","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.title","nameWithType":"SceneCollectionTemplate.title"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection*","name":"CreateCollection","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateCollection_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateCollection","nameWithType":"SceneCollectionTemplate.CreateCollection"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.Apply*","name":"Apply","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_Apply_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.Apply","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.Apply","nameWithType":"SceneCollectionTemplate.Apply"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder*","name":"CreateTemplateInCurrentFolder","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateTemplateInCurrentFolder_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplateInCurrentFolder","nameWithType":"SceneCollectionTemplate.CreateTemplateInCurrentFolder"},{"uid":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate*","name":"CreateTemplate","href":"~/api/AdvancedSceneManager.Models.SceneCollectionTemplate.yml#AdvancedSceneManager_Models_SceneCollectionTemplate_CreateTemplate_","commentId":"Overload:AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneCollectionTemplate.CreateTemplate","nameWithType":"SceneCollectionTemplate.CreateTemplate"}],"api/AdvancedSceneManager.Models.SceneOpenBehavior.yml":[{"uid":"AdvancedSceneManager.Models.SceneOpenBehavior","name":"SceneOpenBehavior","href":"~/api/AdvancedSceneManager.Models.SceneOpenBehavior.yml","commentId":"T:AdvancedSceneManager.Models.SceneOpenBehavior","fullName":"AdvancedSceneManager.Models.SceneOpenBehavior","nameWithType":"SceneOpenBehavior"},{"uid":"AdvancedSceneManager.Models.SceneOpenBehavior.OpenNormally","name":"OpenNormally","href":"~/api/AdvancedSceneManager.Models.SceneOpenBehavior.yml#AdvancedSceneManager_Models_SceneOpenBehavior_OpenNormally","commentId":"F:AdvancedSceneManager.Models.SceneOpenBehavior.OpenNormally","fullName":"AdvancedSceneManager.Models.SceneOpenBehavior.OpenNormally","nameWithType":"SceneOpenBehavior.OpenNormally"},{"uid":"AdvancedSceneManager.Models.SceneOpenBehavior.DoNotOpenInCollection","name":"DoNotOpenInCollection","href":"~/api/AdvancedSceneManager.Models.SceneOpenBehavior.yml#AdvancedSceneManager_Models_SceneOpenBehavior_DoNotOpenInCollection","commentId":"F:AdvancedSceneManager.Models.SceneOpenBehavior.DoNotOpenInCollection","fullName":"AdvancedSceneManager.Models.SceneOpenBehavior.DoNotOpenInCollection","nameWithType":"SceneOpenBehavior.DoNotOpenInCollection"}],"api/AdvancedSceneManager.Utility.DictionaryUtility.yml":[{"uid":"AdvancedSceneManager.Utility.DictionaryUtility","name":"DictionaryUtility","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml","commentId":"T:AdvancedSceneManager.Utility.DictionaryUtility","fullName":"AdvancedSceneManager.Utility.DictionaryUtility","nameWithType":"DictionaryUtility"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey``2(System.Collections.Generic.Dictionary{``0,``1},``0)","name":"WithNullKey<TKey, TValue>(Dictionary<TKey, TValue>, TKey)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_WithNullKey__2_System_Collections_Generic_Dictionary___0___1____0_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey``2(System.Collections.Generic.Dictionary{``0,``1},``0)","name.vb":"WithNullKey(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey<TKey, TValue>(System.Collections.Generic.Dictionary<TKey, TValue>, TKey)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey(Of TKey, TValue)(System.Collections.Generic.Dictionary(Of TKey, TValue), TKey)","nameWithType":"DictionaryUtility.WithNullKey<TKey, TValue>(Dictionary<TKey, TValue>, TKey)","nameWithType.vb":"DictionaryUtility.WithNullKey(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Set``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name":"Set<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Set__2_System_Collections_Generic_Dictionary___0___1____0___1_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.Set``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name.vb":"Set(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Set<TKey, TValue>(System.Collections.Generic.Dictionary<TKey, TValue>, TKey, TValue)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.Set(Of TKey, TValue)(System.Collections.Generic.Dictionary(Of TKey, TValue), TKey, TValue)","nameWithType":"DictionaryUtility.Set<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","nameWithType.vb":"DictionaryUtility.Set(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded``2(System.Collections.Generic.Dictionary{``0,``1},``0)","name":"EnsureAdded<TKey, TValue>(Dictionary<TKey, TValue>, TKey)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_EnsureAdded__2_System_Collections_Generic_Dictionary___0___1____0_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded``2(System.Collections.Generic.Dictionary{``0,``1},``0)","name.vb":"EnsureAdded(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded<TKey, TValue>(System.Collections.Generic.Dictionary<TKey, TValue>, TKey)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded(Of TKey, TValue)(System.Collections.Generic.Dictionary(Of TKey, TValue), TKey)","nameWithType":"DictionaryUtility.EnsureAdded<TKey, TValue>(Dictionary<TKey, TValue>, TKey)","nameWithType.vb":"DictionaryUtility.EnsureAdded(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Add``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name":"Add<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Add__2_System_Collections_Generic_Dictionary___0___1____0___1_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.Add``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name.vb":"Add(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Add<TKey, TValue>(System.Collections.Generic.Dictionary<TKey, TValue>, TKey, TValue)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.Add(Of TKey, TValue)(System.Collections.Generic.Dictionary(Of TKey, TValue), TKey, TValue)","nameWithType":"DictionaryUtility.Add<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","nameWithType.vb":"DictionaryUtility.Add(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Add``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2)","name":"Add<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Add__3_System_Collections_Generic_Dictionary___0___1____0___2_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.Add``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2)","name.vb":"Add(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Add<TKey, TList, TItem>(System.Collections.Generic.Dictionary<TKey, TList>, TKey, TItem)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.Add(Of TKey, TList, TItem)(System.Collections.Generic.Dictionary(Of TKey, TList), TKey, TItem)","nameWithType":"DictionaryUtility.Add<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem)","nameWithType.vb":"DictionaryUtility.Add(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange``3(System.Collections.Generic.Dictionary{``0,``1},``0,System.Collections.Generic.IEnumerable{``2})","name":"AddRange<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, IEnumerable<TItem>)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_AddRange__3_System_Collections_Generic_Dictionary___0___1____0_System_Collections_Generic_IEnumerable___2__","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.AddRange``3(System.Collections.Generic.Dictionary{``0,``1},``0,System.Collections.Generic.IEnumerable{``2})","name.vb":"AddRange(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, IEnumerable(Of TItem))","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange<TKey, TList, TItem>(System.Collections.Generic.Dictionary<TKey, TList>, TKey, System.Collections.Generic.IEnumerable<TItem>)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange(Of TKey, TList, TItem)(System.Collections.Generic.Dictionary(Of TKey, TList), TKey, System.Collections.Generic.IEnumerable(Of TItem))","nameWithType":"DictionaryUtility.AddRange<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, IEnumerable<TItem>)","nameWithType.vb":"DictionaryUtility.AddRange(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, IEnumerable(Of TItem))"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2[])","name":"AddRange<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem[])","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_AddRange__3_System_Collections_Generic_Dictionary___0___1____0___2___","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.AddRange``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2[])","name.vb":"AddRange(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem())","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange<TKey, TList, TItem>(System.Collections.Generic.Dictionary<TKey, TList>, TKey, TItem[])","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange(Of TKey, TList, TItem)(System.Collections.Generic.Dictionary(Of TKey, TList), TKey, TItem())","nameWithType":"DictionaryUtility.AddRange<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem[])","nameWithType.vb":"DictionaryUtility.AddRange(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem())"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Remove``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2)","name":"Remove<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Remove__3_System_Collections_Generic_Dictionary___0___1____0___2_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.Remove``3(System.Collections.Generic.Dictionary{``0,``1},``0,``2)","name.vb":"Remove(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Remove<TKey, TList, TItem>(System.Collections.Generic.Dictionary<TKey, TList>, TKey, TItem)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.Remove(Of TKey, TList, TItem)(System.Collections.Generic.Dictionary(Of TKey, TList), TKey, TItem)","nameWithType":"DictionaryUtility.Remove<TKey, TList, TItem>(Dictionary<TKey, TList>, TKey, TItem)","nameWithType.vb":"DictionaryUtility.Remove(Of TKey, TList, TItem)(Dictionary(Of TKey, TList), TKey, TItem)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.GetValue``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name":"GetValue<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_GetValue__2_System_Collections_Generic_Dictionary___0___1____0___1_","commentId":"M:AdvancedSceneManager.Utility.DictionaryUtility.GetValue``2(System.Collections.Generic.Dictionary{``0,``1},``0,``1)","name.vb":"GetValue(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.GetValue<TKey, TValue>(System.Collections.Generic.Dictionary<TKey, TValue>, TKey, TValue)","fullName.vb":"AdvancedSceneManager.Utility.DictionaryUtility.GetValue(Of TKey, TValue)(System.Collections.Generic.Dictionary(Of TKey, TValue), TKey, TValue)","nameWithType":"DictionaryUtility.GetValue<TKey, TValue>(Dictionary<TKey, TValue>, TKey, TValue)","nameWithType.vb":"DictionaryUtility.GetValue(Of TKey, TValue)(Dictionary(Of TKey, TValue), TKey, TValue)"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey*","name":"WithNullKey","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_WithNullKey_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.WithNullKey","nameWithType":"DictionaryUtility.WithNullKey"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Set*","name":"Set","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Set_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.Set","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Set","nameWithType":"DictionaryUtility.Set"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded*","name":"EnsureAdded","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_EnsureAdded_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.EnsureAdded","nameWithType":"DictionaryUtility.EnsureAdded"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Add*","name":"Add","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Add_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.Add","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Add","nameWithType":"DictionaryUtility.Add"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange*","name":"AddRange","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_AddRange_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.AddRange","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.AddRange","nameWithType":"DictionaryUtility.AddRange"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_Remove_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.Remove","nameWithType":"DictionaryUtility.Remove"},{"uid":"AdvancedSceneManager.Utility.DictionaryUtility.GetValue*","name":"GetValue","href":"~/api/AdvancedSceneManager.Utility.DictionaryUtility.yml#AdvancedSceneManager_Utility_DictionaryUtility_GetValue_","commentId":"Overload:AdvancedSceneManager.Utility.DictionaryUtility.GetValue","isSpec":"True","fullName":"AdvancedSceneManager.Utility.DictionaryUtility.GetValue","nameWithType":"DictionaryUtility.GetValue"}],"api/AdvancedSceneManager.Utility.GuidReference.Editor.yml":[{"uid":"AdvancedSceneManager.Utility.GuidReference.Editor","name":"GuidReference.Editor","href":"~/api/AdvancedSceneManager.Utility.GuidReference.Editor.yml","commentId":"T:AdvancedSceneManager.Utility.GuidReference.Editor","fullName":"AdvancedSceneManager.Utility.GuidReference.Editor","nameWithType":"GuidReference.Editor"},{"uid":"AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI","name":"OnInspectorGUI()","href":"~/api/AdvancedSceneManager.Utility.GuidReference.Editor.yml#AdvancedSceneManager_Utility_GuidReference_Editor_OnInspectorGUI","commentId":"M:AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI","fullName":"AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI()","nameWithType":"GuidReference.Editor.OnInspectorGUI()"},{"uid":"AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins","name":"UseDefaultMargins()","href":"~/api/AdvancedSceneManager.Utility.GuidReference.Editor.yml#AdvancedSceneManager_Utility_GuidReference_Editor_UseDefaultMargins","commentId":"M:AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins","fullName":"AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins()","nameWithType":"GuidReference.Editor.UseDefaultMargins()"},{"uid":"AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI*","name":"OnInspectorGUI","href":"~/api/AdvancedSceneManager.Utility.GuidReference.Editor.yml#AdvancedSceneManager_Utility_GuidReference_Editor_OnInspectorGUI_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReference.Editor.OnInspectorGUI","nameWithType":"GuidReference.Editor.OnInspectorGUI"},{"uid":"AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins*","name":"UseDefaultMargins","href":"~/api/AdvancedSceneManager.Utility.GuidReference.Editor.yml#AdvancedSceneManager_Utility_GuidReference_Editor_UseDefaultMargins_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReference.Editor.UseDefaultMargins","nameWithType":"GuidReference.Editor.UseDefaultMargins"}],"api/AdvancedSceneManager.Utility.yml":[{"uid":"AdvancedSceneManager.Utility","name":"AdvancedSceneManager.Utility","href":"~/api/AdvancedSceneManager.Utility.yml","commentId":"N:AdvancedSceneManager.Utility","fullName":"AdvancedSceneManager.Utility","nameWithType":"AdvancedSceneManager.Utility"}],"api/AdvancedSceneManager.yml":[{"uid":"AdvancedSceneManager","name":"AdvancedSceneManager","href":"~/api/AdvancedSceneManager.yml","commentId":"N:AdvancedSceneManager","fullName":"AdvancedSceneManager","nameWithType":"AdvancedSceneManager"}],"api/AdvancedSceneManager.Callbacks.CombineNull.yml":[{"uid":"AdvancedSceneManager.Callbacks.CombineNull","name":"CombineNull","href":"~/api/AdvancedSceneManager.Callbacks.CombineNull.yml","commentId":"T:AdvancedSceneManager.Callbacks.CombineNull","fullName":"AdvancedSceneManager.Callbacks.CombineNull","nameWithType":"CombineNull"},{"uid":"AdvancedSceneManager.Callbacks.CombineNull.value","name":"value","href":"~/api/AdvancedSceneManager.Callbacks.CombineNull.yml#AdvancedSceneManager_Callbacks_CombineNull_value","commentId":"F:AdvancedSceneManager.Callbacks.CombineNull.value","fullName":"AdvancedSceneManager.Callbacks.CombineNull.value","nameWithType":"CombineNull.value"},{"uid":"AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull(AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","name":"IsCombineNull(CoroutineDiagHelper.SubroutineDetails)","href":"~/api/AdvancedSceneManager.Callbacks.CombineNull.yml#AdvancedSceneManager_Callbacks_CombineNull_IsCombineNull_AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SubroutineDetails_","commentId":"M:AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull(AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","fullName":"AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull(AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SubroutineDetails)","nameWithType":"CombineNull.IsCombineNull(CoroutineDiagHelper.SubroutineDetails)"},{"uid":"AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull*","name":"IsCombineNull","href":"~/api/AdvancedSceneManager.Callbacks.CombineNull.yml#AdvancedSceneManager_Callbacks_CombineNull_IsCombineNull_","commentId":"Overload:AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CombineNull.IsCombineNull","nameWithType":"CombineNull.IsCombineNull"}],"api/AdvancedSceneManager.Callbacks.ISceneManagerCallbackBase.yml":[{"uid":"AdvancedSceneManager.Callbacks.ISceneManagerCallbackBase","name":"ISceneManagerCallbackBase","href":"~/api/AdvancedSceneManager.Callbacks.ISceneManagerCallbackBase.yml","commentId":"T:AdvancedSceneManager.Callbacks.ISceneManagerCallbackBase","fullName":"AdvancedSceneManager.Callbacks.ISceneManagerCallbackBase","nameWithType":"ISceneManagerCallbackBase"}],"api/AdvancedSceneManager.Callbacks.Serializable-2.yml":[{"uid":"AdvancedSceneManager.Callbacks.Serializable`2","name":"Serializable<T, TValue>","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml","commentId":"T:AdvancedSceneManager.Callbacks.Serializable`2","name.vb":"Serializable(Of T, TValue)","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue)","nameWithType":"Serializable<T, TValue>","nameWithType.vb":"Serializable(Of T, TValue)"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.value","name":"value","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_value","commentId":"P:AdvancedSceneManager.Callbacks.Serializable`2.value","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.value","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).value","nameWithType":"Serializable<T, TValue>.value","nameWithType.vb":"Serializable(Of T, TValue).value"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.Convert(`0)","name":"Convert(T)","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_Convert__0_","commentId":"M:AdvancedSceneManager.Callbacks.Serializable`2.Convert(`0)","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.Convert(T)","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).Convert(T)","nameWithType":"Serializable<T, TValue>.Convert(T)","nameWithType.vb":"Serializable(Of T, TValue).Convert(T)"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.ConvertBack(`1)","name":"ConvertBack(TValue)","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_ConvertBack__1_","commentId":"M:AdvancedSceneManager.Callbacks.Serializable`2.ConvertBack(`1)","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.ConvertBack(TValue)","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).ConvertBack(TValue)","nameWithType":"Serializable<T, TValue>.ConvertBack(TValue)","nameWithType.vb":"Serializable(Of T, TValue).ConvertBack(TValue)"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.OnAfterDeserialize","name":"OnAfterDeserialize()","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_OnAfterDeserialize","commentId":"M:AdvancedSceneManager.Callbacks.Serializable`2.OnAfterDeserialize","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.OnAfterDeserialize()","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).OnAfterDeserialize()","nameWithType":"Serializable<T, TValue>.OnAfterDeserialize()","nameWithType.vb":"Serializable(Of T, TValue).OnAfterDeserialize()"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.OnBeforeSerialize","name":"OnBeforeSerialize()","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_OnBeforeSerialize","commentId":"M:AdvancedSceneManager.Callbacks.Serializable`2.OnBeforeSerialize","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.OnBeforeSerialize()","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).OnBeforeSerialize()","nameWithType":"Serializable<T, TValue>.OnBeforeSerialize()","nameWithType.vb":"Serializable(Of T, TValue).OnBeforeSerialize()"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.value*","name":"value","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_value_","commentId":"Overload:AdvancedSceneManager.Callbacks.Serializable`2.value","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.value","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).value","nameWithType":"Serializable<T, TValue>.value","nameWithType.vb":"Serializable(Of T, TValue).value"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.Convert*","name":"Convert","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_Convert_","commentId":"Overload:AdvancedSceneManager.Callbacks.Serializable`2.Convert","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.Convert","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).Convert","nameWithType":"Serializable<T, TValue>.Convert","nameWithType.vb":"Serializable(Of T, TValue).Convert"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.ConvertBack*","name":"ConvertBack","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_ConvertBack_","commentId":"Overload:AdvancedSceneManager.Callbacks.Serializable`2.ConvertBack","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.ConvertBack","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).ConvertBack","nameWithType":"Serializable<T, TValue>.ConvertBack","nameWithType.vb":"Serializable(Of T, TValue).ConvertBack"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.OnAfterDeserialize*","name":"OnAfterDeserialize","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_OnAfterDeserialize_","commentId":"Overload:AdvancedSceneManager.Callbacks.Serializable`2.OnAfterDeserialize","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.OnAfterDeserialize","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).OnAfterDeserialize","nameWithType":"Serializable<T, TValue>.OnAfterDeserialize","nameWithType.vb":"Serializable(Of T, TValue).OnAfterDeserialize"},{"uid":"AdvancedSceneManager.Callbacks.Serializable`2.OnBeforeSerialize*","name":"OnBeforeSerialize","href":"~/api/AdvancedSceneManager.Callbacks.Serializable-2.yml#AdvancedSceneManager_Callbacks_Serializable_2_OnBeforeSerialize_","commentId":"Overload:AdvancedSceneManager.Callbacks.Serializable`2.OnBeforeSerialize","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.Serializable<T, TValue>.OnBeforeSerialize","fullName.vb":"AdvancedSceneManager.Callbacks.Serializable(Of T, TValue).OnBeforeSerialize","nameWithType":"Serializable<T, TValue>.OnBeforeSerialize","nameWithType.vb":"Serializable(Of T, TValue).OnBeforeSerialize"}],"api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction","name":"CloseAllUnityScenesAction","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction","nameWithType":"CloseAllUnityScenesAction"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress","nameWithType":"CloseAllUnityScenesAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor","name":"CloseAllUnityScenesAction()","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction__ctor","commentId":"M:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.CloseAllUnityScenesAction()","nameWithType":"CloseAllUnityScenesAction.CloseAllUnityScenesAction()"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor(System.Func{UnityEngine.SceneManagement.Scene})","name":"CloseAllUnityScenesAction(Func<Scene>)","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction__ctor_System_Func_UnityEngine_SceneManagement_Scene__","commentId":"M:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor(System.Func{UnityEngine.SceneManagement.Scene})","name.vb":"CloseAllUnityScenesAction(Func(Of Scene))","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.CloseAllUnityScenesAction(System.Func<UnityEngine.SceneManagement.Scene>)","fullName.vb":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.CloseAllUnityScenesAction(System.Func(Of UnityEngine.SceneManagement.Scene))","nameWithType":"CloseAllUnityScenesAction.CloseAllUnityScenesAction(Func<Scene>)","nameWithType.vb":"CloseAllUnityScenesAction.CloseAllUnityScenesAction(Func(Of Scene))"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"CloseAllUnityScenesAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.reportsProgress","nameWithType":"CloseAllUnityScenesAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor*","name":"CloseAllUnityScenesAction","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.CloseAllUnityScenesAction","nameWithType":"CloseAllUnityScenesAction.CloseAllUnityScenesAction"},{"uid":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.yml#AdvancedSceneManager_Core_Actions_CloseAllUnityScenesAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.CloseAllUnityScenesAction.DoAction","nameWithType":"CloseAllUnityScenesAction.DoAction"}],"api/AdvancedSceneManager.Core.Actions.QuitAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.QuitAction","name":"QuitAction","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.QuitAction","fullName":"AdvancedSceneManager.Core.Actions.QuitAction","nameWithType":"QuitAction"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_reportsProgress","commentId":"P:AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress","nameWithType":"QuitAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit","name":"CancelQuit()","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_CancelQuit","commentId":"M:AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit()","nameWithType":"QuitAction.CancelQuit()"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.isQuitting","name":"isQuitting","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_isQuitting","commentId":"P:AdvancedSceneManager.Core.Actions.QuitAction.isQuitting","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.isQuitting","nameWithType":"QuitAction.isQuitting"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.#ctor(System.Boolean,System.Nullable{UnityEngine.Color},System.Single,System.Boolean,System.Boolean)","name":"QuitAction(Boolean, Nullable<Color>, Single, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction__ctor_System_Boolean_System_Nullable_UnityEngine_Color__System_Single_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Actions.QuitAction.#ctor(System.Boolean,System.Nullable{UnityEngine.Color},System.Single,System.Boolean,System.Boolean)","name.vb":"QuitAction(Boolean, Nullable(Of Color), Single, Boolean, Boolean)","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.QuitAction(System.Boolean, System.Nullable<UnityEngine.Color>, System.Single, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.QuitAction.QuitAction(System.Boolean, System.Nullable(Of UnityEngine.Color), System.Single, System.Boolean, System.Boolean)","nameWithType":"QuitAction.QuitAction(Boolean, Nullable<Color>, Single, Boolean, Boolean)","nameWithType.vb":"QuitAction.QuitAction(Boolean, Nullable(Of Color), Single, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.QuitAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"QuitAction.DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress*","name":"reportsProgress","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_reportsProgress_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.reportsProgress","nameWithType":"QuitAction.reportsProgress"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit*","name":"CancelQuit","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_CancelQuit_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.CancelQuit","nameWithType":"QuitAction.CancelQuit"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.isQuitting*","name":"isQuitting","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_isQuitting_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuitAction.isQuitting","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.isQuitting","nameWithType":"QuitAction.isQuitting"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.#ctor*","name":"QuitAction","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuitAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.QuitAction","nameWithType":"QuitAction.QuitAction"},{"uid":"AdvancedSceneManager.Core.Actions.QuitAction.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.QuitAction.yml#AdvancedSceneManager_Core_Actions_QuitAction_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.QuitAction.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.QuitAction.DoAction","nameWithType":"QuitAction.DoAction"}],"api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI","name":"HierarchyGUIUtility.HierarchyGameObjectGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI","fullName":"AdvancedSceneManager.Editor.Utility.HierarchyGUIUtility.HierarchyGameObjectGUI","nameWithType":"HierarchyGUIUtility.HierarchyGameObjectGUI"}],"api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption","name":"PersistentSceneInEditorUtility.OpenInEditorOption","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorOption"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.Never","name":"Never","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorOption_Never","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.Never","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.Never","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorOption.Never"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.AnySceneOpens","name":"AnySceneOpens","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorOption_AnySceneOpens","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.AnySceneOpens","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.AnySceneOpens","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorOption.AnySceneOpens"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnyOfTheFollowingScenesOpen","name":"WhenAnyOfTheFollowingScenesOpen","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorOption_WhenAnyOfTheFollowingScenesOpen","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnyOfTheFollowingScenesOpen","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnyOfTheFollowingScenesOpen","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnyOfTheFollowingScenesOpen"},{"uid":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnySceneOpensExcept","name":"WhenAnySceneOpensExcept","href":"~/api/AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.yml#AdvancedSceneManager_Editor_Utility_PersistentSceneInEditorUtility_OpenInEditorOption_WhenAnySceneOpensExcept","commentId":"F:AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnySceneOpensExcept","fullName":"AdvancedSceneManager.Editor.Utility.PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnySceneOpensExcept","nameWithType":"PersistentSceneInEditorUtility.OpenInEditorOption.WhenAnySceneOpensExcept"}],"api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion","name":"PromptVersion","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PromptVersion","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion","nameWithType":"PromptVersion"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_title","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptVersion.title","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.title","nameWithType":"PromptVersion.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.Validate(System.String)","name":"Validate(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_Validate_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptVersion.Validate(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.Validate(System.String)","nameWithType":"PromptVersion.Validate(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI(System.String@)","name":"OnContentGUI(ref String)","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_OnContentGUI_System_String__","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI(System.String@)","name.vb":"OnContentGUI(ByRef String)","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI(ref System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI(ByRef System.String)","nameWithType":"PromptVersion.OnContentGUI(ref String)","nameWithType.vb":"PromptVersion.OnContentGUI(ByRef String)"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptVersion.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.title","nameWithType":"PromptVersion.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.Validate*","name":"Validate","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_Validate_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptVersion.Validate","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.Validate","nameWithType":"PromptVersion.Validate"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptVersion.yml#AdvancedSceneManager_Editor_Utility_PromptVersion_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptVersion.OnContentGUI","nameWithType":"PromptVersion.OnContentGUI"}],"api/AdvancedSceneManager.Editor.yml":[{"uid":"AdvancedSceneManager.Editor","name":"AdvancedSceneManager.Editor","href":"~/api/AdvancedSceneManager.Editor.yml","commentId":"N:AdvancedSceneManager.Editor","fullName":"AdvancedSceneManager.Editor","nameWithType":"AdvancedSceneManager.Editor"}],"api/AdvancedSceneManager.Exceptions.CloseSceneException.yml":[{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException","name":"CloseSceneException","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml","commentId":"T:AdvancedSceneManager.Exceptions.CloseSceneException","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException","nameWithType":"CloseSceneException"},{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException.#ctor(AdvancedSceneManager.Models.Scene,UnityEngine.SceneManagement.Scene,AdvancedSceneManager.Models.SceneCollection,System.String)","name":"CloseSceneException(Scene, Scene, SceneCollection, String)","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml#AdvancedSceneManager_Exceptions_CloseSceneException__ctor_AdvancedSceneManager_Models_Scene_UnityEngine_SceneManagement_Scene_AdvancedSceneManager_Models_SceneCollection_System_String_","commentId":"M:AdvancedSceneManager.Exceptions.CloseSceneException.#ctor(AdvancedSceneManager.Models.Scene,UnityEngine.SceneManagement.Scene,AdvancedSceneManager.Models.SceneCollection,System.String)","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException.CloseSceneException(AdvancedSceneManager.Models.Scene, UnityEngine.SceneManagement.Scene, AdvancedSceneManager.Models.SceneCollection, System.String)","nameWithType":"CloseSceneException.CloseSceneException(Scene, Scene, SceneCollection, String)"},{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException.scene","name":"scene","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml#AdvancedSceneManager_Exceptions_CloseSceneException_scene","commentId":"F:AdvancedSceneManager.Exceptions.CloseSceneException.scene","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException.scene","nameWithType":"CloseSceneException.scene"},{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException.unityScene","name":"unityScene","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml#AdvancedSceneManager_Exceptions_CloseSceneException_unityScene","commentId":"F:AdvancedSceneManager.Exceptions.CloseSceneException.unityScene","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException.unityScene","nameWithType":"CloseSceneException.unityScene"},{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException.collection","name":"collection","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml#AdvancedSceneManager_Exceptions_CloseSceneException_collection","commentId":"F:AdvancedSceneManager.Exceptions.CloseSceneException.collection","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException.collection","nameWithType":"CloseSceneException.collection"},{"uid":"AdvancedSceneManager.Exceptions.CloseSceneException.#ctor*","name":"CloseSceneException","href":"~/api/AdvancedSceneManager.Exceptions.CloseSceneException.yml#AdvancedSceneManager_Exceptions_CloseSceneException__ctor_","commentId":"Overload:AdvancedSceneManager.Exceptions.CloseSceneException.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Exceptions.CloseSceneException.CloseSceneException","nameWithType":"CloseSceneException.CloseSceneException"}],"api/AdvancedSceneManager.Models.DynamicCollection.yml":[{"uid":"AdvancedSceneManager.Models.DynamicCollection","name":"DynamicCollection","href":"~/api/AdvancedSceneManager.Models.DynamicCollection.yml","commentId":"T:AdvancedSceneManager.Models.DynamicCollection","fullName":"AdvancedSceneManager.Models.DynamicCollection","nameWithType":"DynamicCollection"},{"uid":"AdvancedSceneManager.Models.DynamicCollection.title","name":"title","href":"~/api/AdvancedSceneManager.Models.DynamicCollection.yml#AdvancedSceneManager_Models_DynamicCollection_title","commentId":"F:AdvancedSceneManager.Models.DynamicCollection.title","fullName":"AdvancedSceneManager.Models.DynamicCollection.title","nameWithType":"DynamicCollection.title"},{"uid":"AdvancedSceneManager.Models.DynamicCollection.isAuto","name":"isAuto","href":"~/api/AdvancedSceneManager.Models.DynamicCollection.yml#AdvancedSceneManager_Models_DynamicCollection_isAuto","commentId":"F:AdvancedSceneManager.Models.DynamicCollection.isAuto","fullName":"AdvancedSceneManager.Models.DynamicCollection.isAuto","nameWithType":"DynamicCollection.isAuto"},{"uid":"AdvancedSceneManager.Models.DynamicCollection.scenes","name":"scenes","href":"~/api/AdvancedSceneManager.Models.DynamicCollection.yml#AdvancedSceneManager_Models_DynamicCollection_scenes","commentId":"F:AdvancedSceneManager.Models.DynamicCollection.scenes","fullName":"AdvancedSceneManager.Models.DynamicCollection.scenes","nameWithType":"DynamicCollection.scenes"}],"api/AdvancedSceneManager.Models.ISceneObject.yml":[{"uid":"AdvancedSceneManager.Models.ISceneObject","name":"ISceneObject","href":"~/api/AdvancedSceneManager.Models.ISceneObject.yml","commentId":"T:AdvancedSceneManager.Models.ISceneObject","fullName":"AdvancedSceneManager.Models.ISceneObject","nameWithType":"ISceneObject"},{"uid":"AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged","name":"OnPropertyChanged()","href":"~/api/AdvancedSceneManager.Models.ISceneObject.yml#AdvancedSceneManager_Models_ISceneObject_OnPropertyChanged","commentId":"M:AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged","fullName":"AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged()","nameWithType":"ISceneObject.OnPropertyChanged()"},{"uid":"AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged*","name":"OnPropertyChanged","href":"~/api/AdvancedSceneManager.Models.ISceneObject.yml#AdvancedSceneManager_Models_ISceneObject_OnPropertyChanged_","commentId":"Overload:AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged","isSpec":"True","fullName":"AdvancedSceneManager.Models.ISceneObject.OnPropertyChanged","nameWithType":"ISceneObject.OnPropertyChanged"}],"api/AdvancedSceneManager.Utility.ASM.yml":[{"uid":"AdvancedSceneManager.Utility.ASM","name":"ASM","href":"~/api/AdvancedSceneManager.Utility.ASM.yml","commentId":"T:AdvancedSceneManager.Utility.ASM","fullName":"AdvancedSceneManager.Utility.ASM","nameWithType":"ASM"},{"uid":"AdvancedSceneManager.Utility.ASM.name","name":"name","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_name","commentId":"P:AdvancedSceneManager.Utility.ASM.name","fullName":"AdvancedSceneManager.Utility.ASM.name","nameWithType":"ASM.name"},{"uid":"AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.SceneCollection)","name":"Open(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Open_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ASM.Open(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.ASM.ReopenCollection","name":"ReopenCollection()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_ReopenCollection","commentId":"M:AdvancedSceneManager.Utility.ASM.ReopenCollection","fullName":"AdvancedSceneManager.Utility.ASM.ReopenCollection()","nameWithType":"ASM.ReopenCollection()"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection(AdvancedSceneManager.Models.SceneCollection)","name":"OpenOrReopenCollection(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenOrReopenCollection_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ASM.OpenOrReopenCollection(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.Scene)","name":"Open(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Open_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.Open(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.Open(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.Reopen(AdvancedSceneManager.Models.Scene)","name":"Reopen(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Reopen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.Reopen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.Reopen(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.Reopen(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenSingle(AdvancedSceneManager.Models.Scene)","name":"OpenSingle(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenSingle_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.OpenSingle(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.OpenSingle(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.OpenSingle(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.Preload(AdvancedSceneManager.Models.Scene)","name":"Preload(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Preload_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.Preload(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.Preload(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.Preload(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.FinishPreload","name":"FinishPreload()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_FinishPreload","commentId":"M:AdvancedSceneManager.Utility.ASM.FinishPreload","fullName":"AdvancedSceneManager.Utility.ASM.FinishPreload()","nameWithType":"ASM.FinishPreload()"},{"uid":"AdvancedSceneManager.Utility.ASM.DiscardPreload","name":"DiscardPreload()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_DiscardPreload","commentId":"M:AdvancedSceneManager.Utility.ASM.DiscardPreload","fullName":"AdvancedSceneManager.Utility.ASM.DiscardPreload()","nameWithType":"ASM.DiscardPreload()"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenOrReopen(AdvancedSceneManager.Models.Scene)","name":"OpenOrReopen(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenOrReopen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.OpenOrReopen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.OpenOrReopen(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.OpenOrReopen(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith(System.String)","name":"OpenWhereNameStartsWith(String)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenWhereNameStartsWith_System_String_","commentId":"M:AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith(System.String)","fullName":"AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith(System.String)","nameWithType":"ASM.OpenWhereNameStartsWith(String)"},{"uid":"AdvancedSceneManager.Utility.ASM.CloseCollection","name":"CloseCollection()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_CloseCollection","commentId":"M:AdvancedSceneManager.Utility.ASM.CloseCollection","fullName":"AdvancedSceneManager.Utility.ASM.CloseCollection()","nameWithType":"ASM.CloseCollection()"},{"uid":"AdvancedSceneManager.Utility.ASM.Close(AdvancedSceneManager.Models.Scene)","name":"Close(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Close_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.Close(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.Close(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.Close(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection)","name":"Toggle(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Toggle_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ASM.Toggle(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"Toggle(SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Toggle_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","fullName":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"ASM.Toggle(SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene)","name":"Toggle(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Toggle_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.Toggle(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene,System.Boolean)","name":"Toggle(Scene, Boolean)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Toggle_AdvancedSceneManager_Models_Scene_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene,System.Boolean)","fullName":"AdvancedSceneManager.Utility.ASM.Toggle(AdvancedSceneManager.Models.Scene, System.Boolean)","nameWithType":"ASM.Toggle(Scene, Boolean)"},{"uid":"AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.SceneCollection)","name":"IsOpen(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_IsOpen_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"ASM.IsOpen(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.Scene)","name":"IsOpen(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_IsOpen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.IsOpen(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.IsOpen(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.SetActiveScene(AdvancedSceneManager.Models.Scene)","name":"SetActiveScene(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_SetActiveScene_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.SetActiveScene(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.SetActiveScene(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.SetActiveScene(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.FindCollections(AdvancedSceneManager.Models.Scene)","name":"FindCollections(Scene)","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_FindCollections_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.ASM.FindCollections(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.ASM.FindCollections(AdvancedSceneManager.Models.Scene)","nameWithType":"ASM.FindCollections(Scene)"},{"uid":"AdvancedSceneManager.Utility.ASM.Quit","name":"Quit()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Quit","commentId":"M:AdvancedSceneManager.Utility.ASM.Quit","fullName":"AdvancedSceneManager.Utility.ASM.Quit()","nameWithType":"ASM.Quit()"},{"uid":"AdvancedSceneManager.Utility.ASM.Restart","name":"Restart()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Restart","commentId":"M:AdvancedSceneManager.Utility.ASM.Restart","fullName":"AdvancedSceneManager.Utility.ASM.Restart()","nameWithType":"ASM.Restart()"},{"uid":"AdvancedSceneManager.Utility.ASM.RestartCollection","name":"RestartCollection()","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_RestartCollection","commentId":"M:AdvancedSceneManager.Utility.ASM.RestartCollection","fullName":"AdvancedSceneManager.Utility.ASM.RestartCollection()","nameWithType":"ASM.RestartCollection()"},{"uid":"AdvancedSceneManager.Utility.ASM.name*","name":"name","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_name_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.name","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.name","nameWithType":"ASM.name"},{"uid":"AdvancedSceneManager.Utility.ASM.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Open_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Open","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Open","nameWithType":"ASM.Open"},{"uid":"AdvancedSceneManager.Utility.ASM.ReopenCollection*","name":"ReopenCollection","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_ReopenCollection_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.ReopenCollection","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.ReopenCollection","nameWithType":"ASM.ReopenCollection"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection*","name":"OpenOrReopenCollection","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenOrReopenCollection_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.OpenOrReopenCollection","nameWithType":"ASM.OpenOrReopenCollection"},{"uid":"AdvancedSceneManager.Utility.ASM.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Reopen_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Reopen","nameWithType":"ASM.Reopen"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenSingle*","name":"OpenSingle","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenSingle_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.OpenSingle","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.OpenSingle","nameWithType":"ASM.OpenSingle"},{"uid":"AdvancedSceneManager.Utility.ASM.Preload*","name":"Preload","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Preload_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Preload","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Preload","nameWithType":"ASM.Preload"},{"uid":"AdvancedSceneManager.Utility.ASM.FinishPreload*","name":"FinishPreload","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_FinishPreload_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.FinishPreload","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.FinishPreload","nameWithType":"ASM.FinishPreload"},{"uid":"AdvancedSceneManager.Utility.ASM.DiscardPreload*","name":"DiscardPreload","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_DiscardPreload_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.DiscardPreload","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.DiscardPreload","nameWithType":"ASM.DiscardPreload"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenOrReopen*","name":"OpenOrReopen","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenOrReopen_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.OpenOrReopen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.OpenOrReopen","nameWithType":"ASM.OpenOrReopen"},{"uid":"AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith*","name":"OpenWhereNameStartsWith","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_OpenWhereNameStartsWith_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.OpenWhereNameStartsWith","nameWithType":"ASM.OpenWhereNameStartsWith"},{"uid":"AdvancedSceneManager.Utility.ASM.CloseCollection*","name":"CloseCollection","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_CloseCollection_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.CloseCollection","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.CloseCollection","nameWithType":"ASM.CloseCollection"},{"uid":"AdvancedSceneManager.Utility.ASM.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Close_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Close","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Close","nameWithType":"ASM.Close"},{"uid":"AdvancedSceneManager.Utility.ASM.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Toggle_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Toggle","nameWithType":"ASM.Toggle"},{"uid":"AdvancedSceneManager.Utility.ASM.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_IsOpen_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.IsOpen","nameWithType":"ASM.IsOpen"},{"uid":"AdvancedSceneManager.Utility.ASM.SetActiveScene*","name":"SetActiveScene","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_SetActiveScene_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.SetActiveScene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.SetActiveScene","nameWithType":"ASM.SetActiveScene"},{"uid":"AdvancedSceneManager.Utility.ASM.FindCollections*","name":"FindCollections","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_FindCollections_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.FindCollections","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.FindCollections","nameWithType":"ASM.FindCollections"},{"uid":"AdvancedSceneManager.Utility.ASM.Quit*","name":"Quit","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Quit_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Quit","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Quit","nameWithType":"ASM.Quit"},{"uid":"AdvancedSceneManager.Utility.ASM.Restart*","name":"Restart","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_Restart_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.Restart","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.Restart","nameWithType":"ASM.Restart"},{"uid":"AdvancedSceneManager.Utility.ASM.RestartCollection*","name":"RestartCollection","href":"~/api/AdvancedSceneManager.Utility.ASM.yml#AdvancedSceneManager_Utility_ASM_RestartCollection_","commentId":"Overload:AdvancedSceneManager.Utility.ASM.RestartCollection","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ASM.RestartCollection","nameWithType":"ASM.RestartCollection"}],"api/AdvancedSceneManager.Utility.CanvasGroupExtensions.yml":[{"uid":"AdvancedSceneManager.Utility.CanvasGroupExtensions","name":"CanvasGroupExtensions","href":"~/api/AdvancedSceneManager.Utility.CanvasGroupExtensions.yml","commentId":"T:AdvancedSceneManager.Utility.CanvasGroupExtensions","fullName":"AdvancedSceneManager.Utility.CanvasGroupExtensions","nameWithType":"CanvasGroupExtensions"},{"uid":"AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade(UnityEngine.CanvasGroup,System.Single,System.Single,System.Boolean)","name":"Fade(CanvasGroup, Single, Single, Boolean)","href":"~/api/AdvancedSceneManager.Utility.CanvasGroupExtensions.yml#AdvancedSceneManager_Utility_CanvasGroupExtensions_Fade_UnityEngine_CanvasGroup_System_Single_System_Single_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade(UnityEngine.CanvasGroup,System.Single,System.Single,System.Boolean)","fullName":"AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade(UnityEngine.CanvasGroup, System.Single, System.Single, System.Boolean)","nameWithType":"CanvasGroupExtensions.Fade(CanvasGroup, Single, Single, Boolean)"},{"uid":"AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade*","name":"Fade","href":"~/api/AdvancedSceneManager.Utility.CanvasGroupExtensions.yml#AdvancedSceneManager_Utility_CanvasGroupExtensions_Fade_","commentId":"Overload:AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade","isSpec":"True","fullName":"AdvancedSceneManager.Utility.CanvasGroupExtensions.Fade","nameWithType":"CanvasGroupExtensions.Fade"}],"api/AdvancedSceneManager.Utility.LerpUtility.yml":[{"uid":"AdvancedSceneManager.Utility.LerpUtility","name":"LerpUtility","href":"~/api/AdvancedSceneManager.Utility.LerpUtility.yml","commentId":"T:AdvancedSceneManager.Utility.LerpUtility","fullName":"AdvancedSceneManager.Utility.LerpUtility","nameWithType":"LerpUtility"},{"uid":"AdvancedSceneManager.Utility.LerpUtility.Lerp(System.Single,System.Single,System.Single,System.Action{System.Single},System.Action)","name":"Lerp(Single, Single, Single, Action<Single>, Action)","href":"~/api/AdvancedSceneManager.Utility.LerpUtility.yml#AdvancedSceneManager_Utility_LerpUtility_Lerp_System_Single_System_Single_System_Single_System_Action_System_Single__System_Action_","commentId":"M:AdvancedSceneManager.Utility.LerpUtility.Lerp(System.Single,System.Single,System.Single,System.Action{System.Single},System.Action)","name.vb":"Lerp(Single, Single, Single, Action(Of Single), Action)","fullName":"AdvancedSceneManager.Utility.LerpUtility.Lerp(System.Single, System.Single, System.Single, System.Action<System.Single>, System.Action)","fullName.vb":"AdvancedSceneManager.Utility.LerpUtility.Lerp(System.Single, System.Single, System.Single, System.Action(Of System.Single), System.Action)","nameWithType":"LerpUtility.Lerp(Single, Single, Single, Action<Single>, Action)","nameWithType.vb":"LerpUtility.Lerp(Single, Single, Single, Action(Of Single), Action)"},{"uid":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector3,UnityEngine.Vector3,System.Single,System.Action{UnityEngine.Vector3},System.Action)","name":"Lerp(Vector3, Vector3, Single, Action<Vector3>, Action)","href":"~/api/AdvancedSceneManager.Utility.LerpUtility.yml#AdvancedSceneManager_Utility_LerpUtility_Lerp_UnityEngine_Vector3_UnityEngine_Vector3_System_Single_System_Action_UnityEngine_Vector3__System_Action_","commentId":"M:AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector3,UnityEngine.Vector3,System.Single,System.Action{UnityEngine.Vector3},System.Action)","name.vb":"Lerp(Vector3, Vector3, Single, Action(Of Vector3), Action)","fullName":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector3, UnityEngine.Vector3, System.Single, System.Action<UnityEngine.Vector3>, System.Action)","fullName.vb":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector3, UnityEngine.Vector3, System.Single, System.Action(Of UnityEngine.Vector3), System.Action)","nameWithType":"LerpUtility.Lerp(Vector3, Vector3, Single, Action<Vector3>, Action)","nameWithType.vb":"LerpUtility.Lerp(Vector3, Vector3, Single, Action(Of Vector3), Action)"},{"uid":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector2,UnityEngine.Vector2,System.Single,System.Action{UnityEngine.Vector2},System.Action)","name":"Lerp(Vector2, Vector2, Single, Action<Vector2>, Action)","href":"~/api/AdvancedSceneManager.Utility.LerpUtility.yml#AdvancedSceneManager_Utility_LerpUtility_Lerp_UnityEngine_Vector2_UnityEngine_Vector2_System_Single_System_Action_UnityEngine_Vector2__System_Action_","commentId":"M:AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector2,UnityEngine.Vector2,System.Single,System.Action{UnityEngine.Vector2},System.Action)","name.vb":"Lerp(Vector2, Vector2, Single, Action(Of Vector2), Action)","fullName":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector2, UnityEngine.Vector2, System.Single, System.Action<UnityEngine.Vector2>, System.Action)","fullName.vb":"AdvancedSceneManager.Utility.LerpUtility.Lerp(UnityEngine.Vector2, UnityEngine.Vector2, System.Single, System.Action(Of UnityEngine.Vector2), System.Action)","nameWithType":"LerpUtility.Lerp(Vector2, Vector2, Single, Action<Vector2>, Action)","nameWithType.vb":"LerpUtility.Lerp(Vector2, Vector2, Single, Action(Of Vector2), Action)"},{"uid":"AdvancedSceneManager.Utility.LerpUtility.Lerp*","name":"Lerp","href":"~/api/AdvancedSceneManager.Utility.LerpUtility.yml#AdvancedSceneManager_Utility_LerpUtility_Lerp_","commentId":"Overload:AdvancedSceneManager.Utility.LerpUtility.Lerp","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LerpUtility.Lerp","nameWithType":"LerpUtility.Lerp"}],"api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml":[{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility","name":"LoadingScreenUtility","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml","commentId":"T:AdvancedSceneManager.Utility.LoadingScreenUtility","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility","nameWithType":"LoadingScreenUtility"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(UnityEngine.SceneManagement.Scene)","name":"IsLoadingScreenOpen(Scene)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsLoadingScreenOpen_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(UnityEngine.SceneManagement.Scene)","nameWithType":"LoadingScreenUtility.IsLoadingScreenOpen(Scene)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Models.Scene)","name":"IsLoadingScreenOpen(Scene)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsLoadingScreenOpen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Models.Scene)","nameWithType":"LoadingScreenUtility.IsLoadingScreenOpen(Scene)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Core.OpenSceneInfo)","name":"IsLoadingScreenOpen(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsLoadingScreenOpen_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"LoadingScreenUtility.IsLoadingScreenOpen(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen","name":"IsAnyLoadingScreenOpen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsAnyLoadingScreenOpen","commentId":"P:AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen","nameWithType":"LoadingScreenUtility.IsAnyLoadingScreenOpen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Single},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name":"OpenLoadingScreen(SceneCollection, Nullable<Single>, Action<LoadingScreen>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_OpenLoadingScreen_AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Single__System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Single},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name.vb":"OpenLoadingScreen(SceneCollection, Nullable(Of Single), Action(Of LoadingScreen))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Single>, System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Single), System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen))","nameWithType":"LoadingScreenUtility.OpenLoadingScreen(SceneCollection, Nullable<Single>, Action<LoadingScreen>)","nameWithType.vb":"LoadingScreenUtility.OpenLoadingScreen(SceneCollection, Nullable(Of Single), Action(Of LoadingScreen))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.Scene,System.Nullable{System.Single},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen},System.String)","name":"OpenLoadingScreen(Scene, Nullable<Single>, Action<LoadingScreen>, String)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_OpenLoadingScreen_AdvancedSceneManager_Models_Scene_System_Nullable_System_Single__System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__System_String_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.Scene,System.Nullable{System.Single},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen},System.String)","name.vb":"OpenLoadingScreen(Scene, Nullable(Of Single), Action(Of LoadingScreen), String)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.Scene, System.Nullable<System.Single>, System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>, System.String)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(AdvancedSceneManager.Models.Scene, System.Nullable(Of System.Single), System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen), System.String)","nameWithType":"LoadingScreenUtility.OpenLoadingScreen(Scene, Nullable<Single>, Action<LoadingScreen>, String)","nameWithType.vb":"LoadingScreenUtility.OpenLoadingScreen(Scene, Nullable(Of Single), Action(Of LoadingScreen), String)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen``1(AdvancedSceneManager.Models.Scene,System.Nullable{System.Single},System.Action{``0},System.String)","name":"OpenLoadingScreen<T>(Scene, Nullable<Single>, Action<T>, String)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_OpenLoadingScreen__1_AdvancedSceneManager_Models_Scene_System_Nullable_System_Single__System_Action___0__System_String_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen``1(AdvancedSceneManager.Models.Scene,System.Nullable{System.Single},System.Action{``0},System.String)","name.vb":"OpenLoadingScreen(Of T)(Scene, Nullable(Of Single), Action(Of T), String)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen<T>(AdvancedSceneManager.Models.Scene, System.Nullable<System.Single>, System.Action<T>, System.String)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen(Of T)(AdvancedSceneManager.Models.Scene, System.Nullable(Of System.Single), System.Action(Of T), System.String)","nameWithType":"LoadingScreenUtility.OpenLoadingScreen<T>(Scene, Nullable<Single>, Action<T>, String)","nameWithType.vb":"LoadingScreenUtility.OpenLoadingScreen(Of T)(Scene, Nullable(Of Single), Action(Of T), String)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Models.Scene)","name":"CloseLoadingScreen(Scene)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_CloseLoadingScreen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Models.Scene)","nameWithType":"LoadingScreenUtility.CloseLoadingScreen(Scene)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Callbacks.LoadingScreen)","name":"CloseLoadingScreen(LoadingScreen)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_CloseLoadingScreen_AdvancedSceneManager_Callbacks_LoadingScreen_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Callbacks.LoadingScreen)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen(AdvancedSceneManager.Callbacks.LoadingScreen)","nameWithType":"LoadingScreenUtility.CloseLoadingScreen(LoadingScreen)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll","name":"CloseAll()","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_CloseAll","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll()","nameWithType":"LoadingScreenUtility.CloseAll()"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen(AdvancedSceneManager.Models.SceneCollection)","name":"FindLoadingScreen(SceneCollection)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FindLoadingScreen_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"LoadingScreenUtility.FindLoadingScreen(SceneCollection)"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.fade","name":"fade","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_fade","commentId":"P:AdvancedSceneManager.Utility.LoadingScreenUtility.fade","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.fade","nameWithType":"LoadingScreenUtility.fade"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Func{System.Collections.IEnumerator},System.Single,System.Nullable{UnityEngine.Color})","name":"DoActionWithFade(Func<IEnumerator>, Single, Nullable<Color>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoActionWithFade_System_Func_System_Collections_IEnumerator__System_Single_System_Nullable_UnityEngine_Color__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Func{System.Collections.IEnumerator},System.Single,System.Nullable{UnityEngine.Color})","name.vb":"DoActionWithFade(Func(Of IEnumerator), Single, Nullable(Of Color))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Func<System.Collections.IEnumerator>, System.Single, System.Nullable<UnityEngine.Color>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Func(Of System.Collections.IEnumerator), System.Single, System.Nullable(Of UnityEngine.Color))","nameWithType":"LoadingScreenUtility.DoActionWithFade(Func<IEnumerator>, Single, Nullable<Color>)","nameWithType.vb":"LoadingScreenUtility.DoActionWithFade(Func(Of IEnumerator), Single, Nullable(Of Color))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Action,System.Single,System.Nullable{UnityEngine.Color})","name":"DoActionWithFade(Action, Single, Nullable<Color>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoActionWithFade_System_Action_System_Single_System_Nullable_UnityEngine_Color__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Action,System.Single,System.Nullable{UnityEngine.Color})","name.vb":"DoActionWithFade(Action, Single, Nullable(Of Color))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Action, System.Single, System.Nullable<UnityEngine.Color>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade(System.Action, System.Single, System.Nullable(Of UnityEngine.Color))","nameWithType":"LoadingScreenUtility.DoActionWithFade(Action, Single, Nullable<Color>)","nameWithType.vb":"LoadingScreenUtility.DoActionWithFade(Action, Single, Nullable(Of Color))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut(System.Single,System.Nullable{UnityEngine.Color})","name":"FadeOut(Single, Nullable<Color>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FadeOut_System_Single_System_Nullable_UnityEngine_Color__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut(System.Single,System.Nullable{UnityEngine.Color})","name.vb":"FadeOut(Single, Nullable(Of Color))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut(System.Single, System.Nullable<UnityEngine.Color>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut(System.Single, System.Nullable(Of UnityEngine.Color))","nameWithType":"LoadingScreenUtility.FadeOut(Single, Nullable<Color>)","nameWithType.vb":"LoadingScreenUtility.FadeOut(Single, Nullable(Of Color))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn(AdvancedSceneManager.Callbacks.LoadingScreen,System.Single,System.Nullable{UnityEngine.Color})","name":"FadeIn(LoadingScreen, Single, Nullable<Color>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FadeIn_AdvancedSceneManager_Callbacks_LoadingScreen_System_Single_System_Nullable_UnityEngine_Color__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn(AdvancedSceneManager.Callbacks.LoadingScreen,System.Single,System.Nullable{UnityEngine.Color})","name.vb":"FadeIn(LoadingScreen, Single, Nullable(Of Color))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn(AdvancedSceneManager.Callbacks.LoadingScreen, System.Single, System.Nullable<UnityEngine.Color>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn(AdvancedSceneManager.Callbacks.LoadingScreen, System.Single, System.Nullable(Of UnityEngine.Color))","nameWithType":"LoadingScreenUtility.FadeIn(LoadingScreen, Single, Nullable<Color>)","nameWithType.vb":"LoadingScreenUtility.FadeIn(LoadingScreen, Single, Nullable(Of Color))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene,System.Action,System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name":"DoAction(Scene, Action, Action<LoadingScreen>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoAction_AdvancedSceneManager_Models_Scene_System_Action_System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene,System.Action,System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name.vb":"DoAction(Scene, Action, Action(Of LoadingScreen))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene, System.Action, System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene, System.Action, System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen))","nameWithType":"LoadingScreenUtility.DoAction(Scene, Action, Action<LoadingScreen>)","nameWithType.vb":"LoadingScreenUtility.DoAction(Scene, Action, Action(Of LoadingScreen))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene,System.Func{System.Collections.IEnumerator},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name":"DoAction(Scene, Func<IEnumerator>, Action<LoadingScreen>)","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoAction_AdvancedSceneManager_Models_Scene_System_Func_System_Collections_IEnumerator__System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__","commentId":"M:AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene,System.Func{System.Collections.IEnumerator},System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name.vb":"DoAction(Scene, Func(Of IEnumerator), Action(Of LoadingScreen))","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene, System.Func<System.Collections.IEnumerator>, System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>)","fullName.vb":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction(AdvancedSceneManager.Models.Scene, System.Func(Of System.Collections.IEnumerator), System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen))","nameWithType":"LoadingScreenUtility.DoAction(Scene, Func<IEnumerator>, Action<LoadingScreen>)","nameWithType.vb":"LoadingScreenUtility.DoAction(Scene, Func(Of IEnumerator), Action(Of LoadingScreen))"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens","name":"loadingScreens","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_loadingScreens","commentId":"P:AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens","nameWithType":"LoadingScreenUtility.loadingScreens"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen*","name":"IsLoadingScreenOpen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsLoadingScreenOpen_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsLoadingScreenOpen","nameWithType":"LoadingScreenUtility.IsLoadingScreenOpen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen*","name":"IsAnyLoadingScreenOpen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_IsAnyLoadingScreenOpen_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.IsAnyLoadingScreenOpen","nameWithType":"LoadingScreenUtility.IsAnyLoadingScreenOpen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen*","name":"OpenLoadingScreen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_OpenLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.OpenLoadingScreen","nameWithType":"LoadingScreenUtility.OpenLoadingScreen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen*","name":"CloseLoadingScreen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_CloseLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseLoadingScreen","nameWithType":"LoadingScreenUtility.CloseLoadingScreen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll*","name":"CloseAll","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_CloseAll_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.CloseAll","nameWithType":"LoadingScreenUtility.CloseAll"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen*","name":"FindLoadingScreen","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FindLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FindLoadingScreen","nameWithType":"LoadingScreenUtility.FindLoadingScreen"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.fade*","name":"fade","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_fade_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.fade","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.fade","nameWithType":"LoadingScreenUtility.fade"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade*","name":"DoActionWithFade","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoActionWithFade_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoActionWithFade","nameWithType":"LoadingScreenUtility.DoActionWithFade"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut*","name":"FadeOut","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FadeOut_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeOut","nameWithType":"LoadingScreenUtility.FadeOut"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn*","name":"FadeIn","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_FadeIn_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.FadeIn","nameWithType":"LoadingScreenUtility.FadeIn"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_DoAction_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.DoAction","nameWithType":"LoadingScreenUtility.DoAction"},{"uid":"AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens*","name":"loadingScreens","href":"~/api/AdvancedSceneManager.Utility.LoadingScreenUtility.yml#AdvancedSceneManager_Utility_LoadingScreenUtility_loadingScreens_","commentId":"Overload:AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens","isSpec":"True","fullName":"AdvancedSceneManager.Utility.LoadingScreenUtility.loadingScreens","nameWithType":"LoadingScreenUtility.loadingScreens"}],"api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml":[{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails","name":"CoroutineDiagHelper.CallerDetails","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml","commentId":"T:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails","nameWithType":"CoroutineDiagHelper.CallerDetails"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.className","name":"className","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_className","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.className","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.className","nameWithType":"CoroutineDiagHelper.CallerDetails.className"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.method","name":"method","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_method","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.method","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.method","nameWithType":"CoroutineDiagHelper.CallerDetails.method"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.methodParameters","name":"methodParameters","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_methodParameters","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.methodParameters","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.methodParameters","nameWithType":"CoroutineDiagHelper.CallerDetails.methodParameters"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.file","name":"file","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_file","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.file","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.file","nameWithType":"CoroutineDiagHelper.CallerDetails.file"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.line","name":"line","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_line","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.line","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.line","nameWithType":"CoroutineDiagHelper.CallerDetails.line"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_ToString","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString()","nameWithType":"CoroutineDiagHelper.CallerDetails.ToString()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_CallerDetails_ToString_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CallerDetails.ToString","nameWithType":"CoroutineDiagHelper.CallerDetails.ToString"}],"api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml":[{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper","name":"CoroutineDiagHelper","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml","commentId":"T:AdvancedSceneManager.Callbacks.CoroutineDiagHelper","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper","nameWithType":"CoroutineDiagHelper"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startTime","name":"startTime","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_startTime","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startTime","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startTime","nameWithType":"CoroutineDiagHelper.startTime"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startFrame","name":"startFrame","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_startFrame","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startFrame","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.startFrame","nameWithType":"CoroutineDiagHelper.startFrame"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.caller","name":"caller","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_caller","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.caller","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.caller","nameWithType":"CoroutineDiagHelper.caller"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isParallel","name":"isParallel","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_isParallel","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isParallel","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isParallel","nameWithType":"CoroutineDiagHelper.isParallel"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel(System.Boolean)","name":"SetParallel(Boolean)","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SetParallel_System_Boolean_","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel(System.Boolean)","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel(System.Boolean)","nameWithType":"CoroutineDiagHelper.SetParallel(Boolean)"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.description","name":"description","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_description","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.description","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.description","nameWithType":"CoroutineDiagHelper.description"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.details","name":"details","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_details","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.details","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.details","nameWithType":"CoroutineDiagHelper.details"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.duration","name":"duration","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_duration","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.duration","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.duration","nameWithType":"CoroutineDiagHelper.duration"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.durationFrames","name":"durationFrames","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_durationFrames","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.durationFrames","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.durationFrames","nameWithType":"CoroutineDiagHelper.durationFrames"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isPaused","name":"isPaused","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_isPaused","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isPaused","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isPaused","nameWithType":"CoroutineDiagHelper.isPaused"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isComplete","name":"isComplete","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_isComplete","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isComplete","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.isComplete","nameWithType":"CoroutineDiagHelper.isComplete"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.wasCancelled","name":"wasCancelled","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_wasCancelled","commentId":"F:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.wasCancelled","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.wasCancelled","nameWithType":"CoroutineDiagHelper.wasCancelled"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor","name":"CoroutineDiagHelper()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper__ctor","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CoroutineDiagHelper()","nameWithType":"CoroutineDiagHelper.CoroutineDiagHelper()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor(System.ValueTuple{System.Reflection.MethodBase,System.String,System.Int32},System.String)","name":"CoroutineDiagHelper((MethodBase method, String file, Int32 line), String)","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper__ctor_System_ValueTuple_System_Reflection_MethodBase_System_String_System_Int32__System_String_","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor(System.ValueTuple{System.Reflection.MethodBase,System.String,System.Int32},System.String)","name.vb":"CoroutineDiagHelper((method As MethodBase, file As String, line As Int32)(Of MethodBase, String, Int32), String)","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CoroutineDiagHelper(System.ValueTuple<System.Reflection.MethodBase, System.String, System.Int32>, System.String)","fullName.vb":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CoroutineDiagHelper(System.ValueTuple(Of System.Reflection.MethodBase, System.String, System.Int32), System.String)","nameWithType":"CoroutineDiagHelper.CoroutineDiagHelper((MethodBase method, String file, Int32 line), String)","nameWithType.vb":"CoroutineDiagHelper.CoroutineDiagHelper((method As MethodBase, file As String, line As Int32)(Of MethodBase, String, Int32), String)"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset","name":"diagOffset","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_diagOffset","commentId":"P:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset","nameWithType":"CoroutineDiagHelper.diagOffset"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor","name":"ViewCallerInCodeEditor()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_ViewCallerInCodeEditor","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor()","nameWithType":"CoroutineDiagHelper.ViewCallerInCodeEditor()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_ToString","commentId":"M:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString()","nameWithType":"CoroutineDiagHelper.ToString()"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel*","name":"SetParallel","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_SetParallel_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.SetParallel","nameWithType":"CoroutineDiagHelper.SetParallel"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor*","name":"CoroutineDiagHelper","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper__ctor_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.CoroutineDiagHelper","nameWithType":"CoroutineDiagHelper.CoroutineDiagHelper"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset*","name":"diagOffset","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_diagOffset_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.diagOffset","nameWithType":"CoroutineDiagHelper.diagOffset"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor*","name":"ViewCallerInCodeEditor","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_ViewCallerInCodeEditor_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ViewCallerInCodeEditor","nameWithType":"CoroutineDiagHelper.ViewCallerInCodeEditor"},{"uid":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Callbacks.CoroutineDiagHelper.yml#AdvancedSceneManager_Callbacks_CoroutineDiagHelper_ToString_","commentId":"Overload:AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.CoroutineDiagHelper.ToString","nameWithType":"CoroutineDiagHelper.ToString"}],"api/AdvancedSceneManager.Callbacks.LoadingScreen.yml":[{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen","name":"LoadingScreen","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml","commentId":"T:AdvancedSceneManager.Callbacks.LoadingScreen","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen","nameWithType":"LoadingScreen"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.onDestroy","name":"onDestroy","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_onDestroy","commentId":"F:AdvancedSceneManager.Callbacks.LoadingScreen.onDestroy","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.onDestroy","nameWithType":"LoadingScreen.onDestroy"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy","name":"OnDestroy()","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnDestroy","commentId":"M:AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy()","nameWithType":"LoadingScreen.OnDestroy()"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.canvas","name":"canvas","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_canvas","commentId":"F:AdvancedSceneManager.Callbacks.LoadingScreen.canvas","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.canvas","nameWithType":"LoadingScreen.canvas"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.operation","name":"operation","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_operation","commentId":"P:AdvancedSceneManager.Callbacks.LoadingScreen.operation","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.operation","nameWithType":"LoadingScreen.operation"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"LoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Callbacks.LoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"LoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged(AdvancedSceneManager.Core.SceneOperation,AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Core.Phase)","name":"OnScenePhaseChanged(SceneOperation, Phase, Phase)","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnScenePhaseChanged_AdvancedSceneManager_Core_SceneOperation_AdvancedSceneManager_Core_Phase_AdvancedSceneManager_Core_Phase_","commentId":"M:AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged(AdvancedSceneManager.Core.SceneOperation,AdvancedSceneManager.Core.Phase,AdvancedSceneManager.Core.Phase)","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged(AdvancedSceneManager.Core.SceneOperation, AdvancedSceneManager.Core.Phase, AdvancedSceneManager.Core.Phase)","nameWithType":"LoadingScreen.OnScenePhaseChanged(SceneOperation, Phase, Phase)"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel(AdvancedSceneManager.Core.SceneOperation)","name":"OnCancel(SceneOperation)","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnCancel_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"LoadingScreen.OnCancel(SceneOperation)"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy*","name":"OnDestroy","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnDestroy_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnDestroy","nameWithType":"LoadingScreen.OnDestroy"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.operation*","name":"operation","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_operation_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.operation","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.operation","nameWithType":"LoadingScreen.operation"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnOpen","nameWithType":"LoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnClose","nameWithType":"LoadingScreen.OnClose"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged*","name":"OnScenePhaseChanged","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnScenePhaseChanged_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnScenePhaseChanged","nameWithType":"LoadingScreen.OnScenePhaseChanged"},{"uid":"AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel*","name":"OnCancel","href":"~/api/AdvancedSceneManager.Callbacks.LoadingScreen.yml#AdvancedSceneManager_Callbacks_LoadingScreen_OnCancel_","commentId":"Overload:AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel","isSpec":"True","fullName":"AdvancedSceneManager.Callbacks.LoadingScreen.OnCancel","nameWithType":"LoadingScreen.OnCancel"}],"api/AdvancedSceneManager.Callbacks.yml":[{"uid":"AdvancedSceneManager.Callbacks","name":"AdvancedSceneManager.Callbacks","href":"~/api/AdvancedSceneManager.Callbacks.yml","commentId":"N:AdvancedSceneManager.Callbacks","fullName":"AdvancedSceneManager.Callbacks","nameWithType":"AdvancedSceneManager.Callbacks"}],"api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml":[{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1","name":"OverridableAction<T>","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml","commentId":"T:AdvancedSceneManager.Core.Actions.OverridableAction`1","name.vb":"OverridableAction(Of T)","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T)","nameWithType":"OverridableAction<T>","nameWithType.vb":"OverridableAction(Of T)"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.overrides","name":"overrides","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_overrides","commentId":"P:AdvancedSceneManager.Core.Actions.OverridableAction`1.overrides","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.overrides","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).overrides","nameWithType":"OverridableAction<T>.overrides","nameWithType.vb":"OverridableAction(Of T).overrides"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.Override(System.String,System.Func{AdvancedSceneManager.Core.SceneManagerBase,`0,System.Collections.IEnumerator})","name":"Override(String, Func<SceneManagerBase, T, IEnumerator>)","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_Override_System_String_System_Func_AdvancedSceneManager_Core_SceneManagerBase__0_System_Collections_IEnumerator__","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.Override(System.String,System.Func{AdvancedSceneManager.Core.SceneManagerBase,`0,System.Collections.IEnumerator})","name.vb":"Override(String, Func(Of SceneManagerBase, T, IEnumerator))","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.Override(System.String, System.Func<AdvancedSceneManager.Core.SceneManagerBase, T, System.Collections.IEnumerator>)","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).Override(System.String, System.Func(Of AdvancedSceneManager.Core.SceneManagerBase, T, System.Collections.IEnumerator))","nameWithType":"OverridableAction<T>.Override(String, Func<SceneManagerBase, T, IEnumerator>)","nameWithType.vb":"OverridableAction(Of T).Override(String, Func(Of SceneManagerBase, T, IEnumerator))"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverride(System.String)","name":"ClearOverride(String)","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ClearOverride_System_String_","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverride(System.String)","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ClearOverride(System.String)","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ClearOverride(System.String)","nameWithType":"OverridableAction<T>.ClearOverride(String)","nameWithType.vb":"OverridableAction(Of T).ClearOverride(String)"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverrides","name":"ClearOverrides()","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ClearOverrides","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverrides","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ClearOverrides()","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ClearOverrides()","nameWithType":"OverridableAction<T>.ClearOverrides()","nameWithType.vb":"OverridableAction(Of T).ClearOverrides()"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_DoAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.DoAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).DoAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"OverridableAction<T>.DoAction(SceneManagerBase)","nameWithType.vb":"OverridableAction(Of T).DoAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","name":"DoNonOverridenAction(SceneManagerBase)","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_DoNonOverridenAction_AdvancedSceneManager_Core_SceneManagerBase_","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).DoNonOverridenAction(AdvancedSceneManager.Core.SceneManagerBase)","nameWithType":"OverridableAction<T>.DoNonOverridenAction(SceneManagerBase)","nameWithType.vb":"OverridableAction(Of T).DoNonOverridenAction(SceneManagerBase)"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.BeforeDoAction(System.Boolean@)","name":"BeforeDoAction(out Boolean)","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_BeforeDoAction_System_Boolean__","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.BeforeDoAction(System.Boolean@)","name.vb":"BeforeDoAction(ByRef Boolean)","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.BeforeDoAction(out System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).BeforeDoAction(ByRef System.Boolean)","nameWithType":"OverridableAction<T>.BeforeDoAction(out Boolean)","nameWithType.vb":"OverridableAction(Of T).BeforeDoAction(ByRef Boolean)"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.lazyScene","name":"lazyScene","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_lazyScene","commentId":"P:AdvancedSceneManager.Core.Actions.OverridableAction`1.lazyScene","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.lazyScene","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).lazyScene","nameWithType":"OverridableAction<T>.lazyScene","nameWithType.vb":"OverridableAction(Of T).lazyScene"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ToString","commentId":"M:AdvancedSceneManager.Core.Actions.OverridableAction`1.ToString","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ToString()","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ToString()","nameWithType":"OverridableAction<T>.ToString()","nameWithType.vb":"OverridableAction(Of T).ToString()"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.overrides*","name":"overrides","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_overrides_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.overrides","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.overrides","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).overrides","nameWithType":"OverridableAction<T>.overrides","nameWithType.vb":"OverridableAction(Of T).overrides"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.Override*","name":"Override","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_Override_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.Override","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.Override","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).Override","nameWithType":"OverridableAction<T>.Override","nameWithType.vb":"OverridableAction(Of T).Override"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverride*","name":"ClearOverride","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ClearOverride_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverride","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ClearOverride","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ClearOverride","nameWithType":"OverridableAction<T>.ClearOverride","nameWithType.vb":"OverridableAction(Of T).ClearOverride"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverrides*","name":"ClearOverrides","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ClearOverrides_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.ClearOverrides","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ClearOverrides","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ClearOverrides","nameWithType":"OverridableAction<T>.ClearOverrides","nameWithType.vb":"OverridableAction(Of T).ClearOverrides"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.DoAction*","name":"DoAction","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_DoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.DoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.DoAction","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).DoAction","nameWithType":"OverridableAction<T>.DoAction","nameWithType.vb":"OverridableAction(Of T).DoAction"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.DoNonOverridenAction*","name":"DoNonOverridenAction","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_DoNonOverridenAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.DoNonOverridenAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.DoNonOverridenAction","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).DoNonOverridenAction","nameWithType":"OverridableAction<T>.DoNonOverridenAction","nameWithType.vb":"OverridableAction(Of T).DoNonOverridenAction"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.BeforeDoAction*","name":"BeforeDoAction","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_BeforeDoAction_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.BeforeDoAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.BeforeDoAction","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).BeforeDoAction","nameWithType":"OverridableAction<T>.BeforeDoAction","nameWithType.vb":"OverridableAction(Of T).BeforeDoAction"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.lazyScene*","name":"lazyScene","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_lazyScene_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.lazyScene","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.lazyScene","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).lazyScene","nameWithType":"OverridableAction<T>.lazyScene","nameWithType.vb":"OverridableAction(Of T).lazyScene"},{"uid":"AdvancedSceneManager.Core.Actions.OverridableAction`1.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Core.Actions.OverridableAction-1.yml#AdvancedSceneManager_Core_Actions_OverridableAction_1_ToString_","commentId":"Overload:AdvancedSceneManager.Core.Actions.OverridableAction`1.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.OverridableAction<T>.ToString","fullName.vb":"AdvancedSceneManager.Core.Actions.OverridableAction(Of T).ToString","nameWithType":"OverridableAction<T>.ToString","nameWithType.vb":"OverridableAction(Of T).ToString"}],"api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseAction","name":"SceneCloseAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneCloseAction","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseAction","nameWithType":"SceneCloseAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","name":"SceneCloseAction(OpenSceneInfo, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseAction__ctor_AdvancedSceneManager_Core_OpenSceneInfo_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseAction.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseAction.SceneCloseAction(AdvancedSceneManager.Core.OpenSceneInfo, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneCloseAction.SceneCloseAction(OpenSceneInfo, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone","name":"OnDone()","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseAction_OnDone","commentId":"M:AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone()","nameWithType":"SceneCloseAction.OnDone()"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseAction.#ctor*","name":"SceneCloseAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneCloseAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseAction.SceneCloseAction","nameWithType":"SceneCloseAction.SceneCloseAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone*","name":"OnDone","href":"~/api/AdvancedSceneManager.Core.Actions.SceneCloseAction.yml#AdvancedSceneManager_Core_Actions_SceneCloseAction_OnDone_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneCloseAction.OnDone","nameWithType":"SceneCloseAction.OnDone"}],"api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml":[{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenAction","name":"SceneOpenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml","commentId":"T:AdvancedSceneManager.Core.Actions.SceneOpenAction","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenAction","nameWithType":"SceneOpenAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenAction.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","name":"SceneOpenAction(Scene, SceneCollection)","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenAction__ctor_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenAction.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenAction.SceneOpenAction(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.SceneCollection)","nameWithType":"SceneOpenAction.SceneOpenAction(Scene, SceneCollection)"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone","name":"OnDone()","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenAction_OnDone","commentId":"M:AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone()","nameWithType":"SceneOpenAction.OnDone()"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenAction.#ctor*","name":"SceneOpenAction","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenAction__ctor_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneOpenAction.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenAction.SceneOpenAction","nameWithType":"SceneOpenAction.SceneOpenAction"},{"uid":"AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone*","name":"OnDone","href":"~/api/AdvancedSceneManager.Core.Actions.SceneOpenAction.yml#AdvancedSceneManager_Core_Actions_SceneOpenAction_OnDone_","commentId":"Overload:AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone","isSpec":"True","fullName":"AdvancedSceneManager.Core.Actions.SceneOpenAction.OnDone","nameWithType":"SceneOpenAction.OnDone"}],"api/AdvancedSceneManager.Core.AssetManagement.yml":[{"uid":"AdvancedSceneManager.Core.AssetManagement","name":"AssetManagement","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml","commentId":"T:AdvancedSceneManager.Core.AssetManagement","fullName":"AdvancedSceneManager.Core.AssetManagement","nameWithType":"AssetManagement"},{"uid":"AdvancedSceneManager.Core.AssetManagement.collections","name":"collections","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_collections","commentId":"P:AdvancedSceneManager.Core.AssetManagement.collections","fullName":"AdvancedSceneManager.Core.AssetManagement.collections","nameWithType":"AssetManagement.collections"},{"uid":"AdvancedSceneManager.Core.AssetManagement.scenes","name":"scenes","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_scenes","commentId":"P:AdvancedSceneManager.Core.AssetManagement.scenes","fullName":"AdvancedSceneManager.Core.AssetManagement.scenes","nameWithType":"AssetManagement.scenes"},{"uid":"AdvancedSceneManager.Core.AssetManagement.profiles","name":"profiles","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_profiles","commentId":"P:AdvancedSceneManager.Core.AssetManagement.profiles","fullName":"AdvancedSceneManager.Core.AssetManagement.profiles","nameWithType":"AssetManagement.profiles"},{"uid":"AdvancedSceneManager.Core.AssetManagement.AssetsChanged","name":"AssetsChanged","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_AssetsChanged","commentId":"E:AdvancedSceneManager.Core.AssetManagement.AssetsChanged","fullName":"AdvancedSceneManager.Core.AssetManagement.AssetsChanged","nameWithType":"AssetManagement.AssetsChanged"},{"uid":"AdvancedSceneManager.Core.AssetManagement.AssetsCleared","name":"AssetsCleared","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_AssetsCleared","commentId":"E:AdvancedSceneManager.Core.AssetManagement.AssetsCleared","fullName":"AdvancedSceneManager.Core.AssetManagement.AssetsCleared","nameWithType":"AssetManagement.AssetsCleared"},{"uid":"AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh","name":"allowAutoRefresh","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_allowAutoRefresh","commentId":"P:AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh","fullName":"AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh","nameWithType":"AssetManagement.allowAutoRefresh"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Rename``1(``0,System.String)","name":"Rename<T>(T, String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Rename__1___0_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Rename``1(``0,System.String)","name.vb":"Rename(Of T)(T, String)","fullName":"AdvancedSceneManager.Core.AssetManagement.Rename<T>(T, System.String)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.Rename(Of T)(T, System.String)","nameWithType":"AssetManagement.Rename<T>(T, String)","nameWithType.vb":"AssetManagement.Rename(Of T)(T, String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Ignore(System.String)","name":"Ignore(String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Ignore_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Ignore(System.String)","fullName":"AdvancedSceneManager.Core.AssetManagement.Ignore(System.String)","nameWithType":"AssetManagement.Ignore(String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.IsIgnored(System.String)","name":"IsIgnored(String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_IsIgnored_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.IsIgnored(System.String)","fullName":"AdvancedSceneManager.Core.AssetManagement.IsIgnored(System.String)","nameWithType":"AssetManagement.IsIgnored(String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindSceneByPath(System.String)","name":"FindSceneByPath(String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindSceneByPath_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.FindSceneByPath(System.String)","fullName":"AdvancedSceneManager.Core.AssetManagement.FindSceneByPath(System.String)","nameWithType":"AssetManagement.FindSceneByPath(String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign","name":"DuplicateProfileAndAssign()","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_DuplicateProfileAndAssign","commentId":"M:AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign","fullName":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign()","nameWithType":"AssetManagement.DuplicateProfileAndAssign()"},{"uid":"AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign(System.Boolean)","name":"CreateProfileAndAssign(Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_CreateProfileAndAssign_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign(System.Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign(System.Boolean)","nameWithType":"AssetManagement.CreateProfileAndAssign(Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfile","name":"DuplicateProfile()","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_DuplicateProfile","commentId":"M:AdvancedSceneManager.Core.AssetManagement.DuplicateProfile","fullName":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfile()","nameWithType":"AssetManagement.DuplicateProfile()"},{"uid":"AdvancedSceneManager.Core.AssetManagement.CreateProfile(System.String,System.Boolean)","name":"CreateProfile(String, Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_CreateProfile_System_String_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.CreateProfile(System.String,System.Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.CreateProfile(System.String, System.Boolean)","nameWithType":"AssetManagement.CreateProfile(String, Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindAssetByID``1(System.String)","name":"FindAssetByID<T>(String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindAssetByID__1_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.FindAssetByID``1(System.String)","name.vb":"FindAssetByID(Of T)(String)","fullName":"AdvancedSceneManager.Core.AssetManagement.FindAssetByID<T>(System.String)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.FindAssetByID(Of T)(System.String)","nameWithType":"AssetManagement.FindAssetByID<T>(String)","nameWithType.vb":"AssetManagement.FindAssetByID(Of T)(String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindAssetByPath``1(System.String)","name":"FindAssetByPath<T>(String)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindAssetByPath__1_System_String_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.FindAssetByPath``1(System.String)","name.vb":"FindAssetByPath(Of T)(String)","fullName":"AdvancedSceneManager.Core.AssetManagement.FindAssetByPath<T>(System.String)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.FindAssetByPath(Of T)(System.String)","nameWithType":"AssetManagement.FindAssetByPath<T>(String)","nameWithType.vb":"AssetManagement.FindAssetByPath(Of T)(String)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Add``1(``0,AdvancedSceneManager.Models.Profile,System.Boolean,System.Boolean)","name":"Add<T>(T, Profile, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Add__1___0_AdvancedSceneManager_Models_Profile_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Add``1(``0,AdvancedSceneManager.Models.Profile,System.Boolean,System.Boolean)","name.vb":"Add(Of T)(T, Profile, Boolean, Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.Add<T>(T, AdvancedSceneManager.Models.Profile, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.Add(Of T)(T, AdvancedSceneManager.Models.Profile, System.Boolean, System.Boolean)","nameWithType":"AssetManagement.Add<T>(T, Profile, Boolean, Boolean)","nameWithType.vb":"AssetManagement.Add(Of T)(T, Profile, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Remove``1(``0)","name":"Remove<T>(T)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Remove__1___0_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Remove``1(``0)","name.vb":"Remove(Of T)(T)","fullName":"AdvancedSceneManager.Core.AssetManagement.Remove<T>(T)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.Remove(Of T)(T)","nameWithType":"AssetManagement.Remove<T>(T)","nameWithType.vb":"AssetManagement.Remove(Of T)(T)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile(AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name":"AddCollectionToProfile(SceneCollection, Profile)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_AddCollectionToProfile_AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile(AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile(AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","nameWithType":"AssetManagement.AddCollectionToProfile(SceneCollection, Profile)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Add(UnityEditor.SceneAsset,System.Boolean)","name":"Add(SceneAsset, Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Add_UnityEditor_SceneAsset_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Add(UnityEditor.SceneAsset,System.Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.Add(UnityEditor.SceneAsset, System.Boolean)","nameWithType":"AssetManagement.Add(SceneAsset, Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Create``1(System.String,System.Action{``0},System.Boolean)","name":"Create<T>(String, Action<T>, Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Create__1_System_String_System_Action___0__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Create``1(System.String,System.Action{``0},System.Boolean)","name.vb":"Create(Of T)(String, Action(Of T), Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.Create<T>(System.String, System.Action<T>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.Create(Of T)(System.String, System.Action(Of T), System.Boolean)","nameWithType":"AssetManagement.Create<T>(String, Action<T>, Boolean)","nameWithType.vb":"AssetManagement.Create(Of T)(String, Action(Of T), Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Create``1(System.String,AdvancedSceneManager.Models.Profile,System.Action{``0},System.Boolean)","name":"Create<T>(String, Profile, Action<T>, Boolean)","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Create__1_System_String_AdvancedSceneManager_Models_Profile_System_Action___0__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Create``1(System.String,AdvancedSceneManager.Models.Profile,System.Action{``0},System.Boolean)","name.vb":"Create(Of T)(String, Profile, Action(Of T), Boolean)","fullName":"AdvancedSceneManager.Core.AssetManagement.Create<T>(System.String, AdvancedSceneManager.Models.Profile, System.Action<T>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.AssetManagement.Create(Of T)(System.String, AdvancedSceneManager.Models.Profile, System.Action(Of T), System.Boolean)","nameWithType":"AssetManagement.Create<T>(String, Profile, Action<T>, Boolean)","nameWithType.vb":"AssetManagement.Create(Of T)(String, Profile, Action(Of T), Boolean)"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Clear","name":"Clear()","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Clear","commentId":"M:AdvancedSceneManager.Core.AssetManagement.Clear","fullName":"AdvancedSceneManager.Core.AssetManagement.Clear()","nameWithType":"AssetManagement.Clear()"},{"uid":"AdvancedSceneManager.Core.AssetManagement.collections*","name":"collections","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_collections_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.collections","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.collections","nameWithType":"AssetManagement.collections"},{"uid":"AdvancedSceneManager.Core.AssetManagement.scenes*","name":"scenes","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_scenes_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.scenes","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.scenes","nameWithType":"AssetManagement.scenes"},{"uid":"AdvancedSceneManager.Core.AssetManagement.profiles*","name":"profiles","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_profiles_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.profiles","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.profiles","nameWithType":"AssetManagement.profiles"},{"uid":"AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh*","name":"allowAutoRefresh","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_allowAutoRefresh_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.allowAutoRefresh","nameWithType":"AssetManagement.allowAutoRefresh"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Rename*","name":"Rename","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Rename_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Rename","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Rename","nameWithType":"AssetManagement.Rename"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Ignore*","name":"Ignore","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Ignore_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Ignore","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Ignore","nameWithType":"AssetManagement.Ignore"},{"uid":"AdvancedSceneManager.Core.AssetManagement.IsIgnored*","name":"IsIgnored","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_IsIgnored_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.IsIgnored","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.IsIgnored","nameWithType":"AssetManagement.IsIgnored"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindSceneByPath*","name":"FindSceneByPath","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindSceneByPath_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.FindSceneByPath","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.FindSceneByPath","nameWithType":"AssetManagement.FindSceneByPath"},{"uid":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign*","name":"DuplicateProfileAndAssign","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_DuplicateProfileAndAssign_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfileAndAssign","nameWithType":"AssetManagement.DuplicateProfileAndAssign"},{"uid":"AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign*","name":"CreateProfileAndAssign","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_CreateProfileAndAssign_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.CreateProfileAndAssign","nameWithType":"AssetManagement.CreateProfileAndAssign"},{"uid":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfile*","name":"DuplicateProfile","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_DuplicateProfile_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.DuplicateProfile","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.DuplicateProfile","nameWithType":"AssetManagement.DuplicateProfile"},{"uid":"AdvancedSceneManager.Core.AssetManagement.CreateProfile*","name":"CreateProfile","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_CreateProfile_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.CreateProfile","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.CreateProfile","nameWithType":"AssetManagement.CreateProfile"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindAssetByID*","name":"FindAssetByID","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindAssetByID_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.FindAssetByID","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.FindAssetByID","nameWithType":"AssetManagement.FindAssetByID"},{"uid":"AdvancedSceneManager.Core.AssetManagement.FindAssetByPath*","name":"FindAssetByPath","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_FindAssetByPath_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.FindAssetByPath","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.FindAssetByPath","nameWithType":"AssetManagement.FindAssetByPath"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Add*","name":"Add","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Add_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Add","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Add","nameWithType":"AssetManagement.Add"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Remove_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Remove","nameWithType":"AssetManagement.Remove"},{"uid":"AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile*","name":"AddCollectionToProfile","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_AddCollectionToProfile_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.AddCollectionToProfile","nameWithType":"AssetManagement.AddCollectionToProfile"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Create*","name":"Create","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Create_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Create","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Create","nameWithType":"AssetManagement.Create"},{"uid":"AdvancedSceneManager.Core.AssetManagement.Clear*","name":"Clear","href":"~/api/AdvancedSceneManager.Core.AssetManagement.yml#AdvancedSceneManager_Core_AssetManagement_Clear_","commentId":"Overload:AdvancedSceneManager.Core.AssetManagement.Clear","isSpec":"True","fullName":"AdvancedSceneManager.Core.AssetManagement.Clear","nameWithType":"AssetManagement.Clear"}],"api/AdvancedSceneManager.Core.Runtime.StartProps.yml":[{"uid":"AdvancedSceneManager.Core.Runtime.StartProps","name":"Runtime.StartProps","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml","commentId":"T:AdvancedSceneManager.Core.Runtime.StartProps","fullName":"AdvancedSceneManager.Core.Runtime.StartProps","nameWithType":"Runtime.StartProps"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.GetDefault","name":"GetDefault()","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_GetDefault","commentId":"M:AdvancedSceneManager.Core.Runtime.StartProps.GetDefault","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.GetDefault()","nameWithType":"Runtime.StartProps.GetDefault()"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.skipSplashScreen","name":"skipSplashScreen","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_skipSplashScreen","commentId":"F:AdvancedSceneManager.Core.Runtime.StartProps.skipSplashScreen","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.skipSplashScreen","nameWithType":"Runtime.StartProps.skipSplashScreen"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.ignoreDoNotOpen","name":"ignoreDoNotOpen","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_ignoreDoNotOpen","commentId":"F:AdvancedSceneManager.Core.Runtime.StartProps.ignoreDoNotOpen","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.ignoreDoNotOpen","nameWithType":"Runtime.StartProps.ignoreDoNotOpen"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.fadeColor","name":"fadeColor","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_fadeColor","commentId":"F:AdvancedSceneManager.Core.Runtime.StartProps.fadeColor","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.fadeColor","nameWithType":"Runtime.StartProps.fadeColor"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.initialFadeDuration","name":"initialFadeDuration","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_initialFadeDuration","commentId":"F:AdvancedSceneManager.Core.Runtime.StartProps.initialFadeDuration","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.initialFadeDuration","nameWithType":"Runtime.StartProps.initialFadeDuration"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.beforeSplashScreenFadeDuration","name":"beforeSplashScreenFadeDuration","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_beforeSplashScreenFadeDuration","commentId":"F:AdvancedSceneManager.Core.Runtime.StartProps.beforeSplashScreenFadeDuration","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.beforeSplashScreenFadeDuration","nameWithType":"Runtime.StartProps.beforeSplashScreenFadeDuration"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection","name":"overrideOpenCollection","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_overrideOpenCollection","commentId":"P:AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection","nameWithType":"Runtime.StartProps.overrideOpenCollection"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.GetDefault*","name":"GetDefault","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_GetDefault_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.StartProps.GetDefault","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.GetDefault","nameWithType":"Runtime.StartProps.GetDefault"},{"uid":"AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection*","name":"overrideOpenCollection","href":"~/api/AdvancedSceneManager.Core.Runtime.StartProps.yml#AdvancedSceneManager_Core_Runtime_StartProps_overrideOpenCollection_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.StartProps.overrideOpenCollection","nameWithType":"Runtime.StartProps.overrideOpenCollection"}],"api/AdvancedSceneManager.Core.Runtime.yml":[{"uid":"AdvancedSceneManager.Core.Runtime","name":"Runtime","href":"~/api/AdvancedSceneManager.Core.Runtime.yml","commentId":"T:AdvancedSceneManager.Core.Runtime","fullName":"AdvancedSceneManager.Core.Runtime","nameWithType":"Runtime"},{"uid":"AdvancedSceneManager.Core.Runtime.isInitialized","name":"isInitialized","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isInitialized","commentId":"P:AdvancedSceneManager.Core.Runtime.isInitialized","fullName":"AdvancedSceneManager.Core.Runtime.isInitialized","nameWithType":"Runtime.isInitialized"},{"uid":"AdvancedSceneManager.Core.Runtime.beforeStart","name":"beforeStart","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_beforeStart","commentId":"E:AdvancedSceneManager.Core.Runtime.beforeStart","fullName":"AdvancedSceneManager.Core.Runtime.beforeStart","nameWithType":"Runtime.beforeStart"},{"uid":"AdvancedSceneManager.Core.Runtime.afterStart","name":"afterStart","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_afterStart","commentId":"E:AdvancedSceneManager.Core.Runtime.afterStart","fullName":"AdvancedSceneManager.Core.Runtime.afterStart","nameWithType":"Runtime.afterStart"},{"uid":"AdvancedSceneManager.Core.Runtime.isBuildMode","name":"isBuildMode","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isBuildMode","commentId":"P:AdvancedSceneManager.Core.Runtime.isBuildMode","fullName":"AdvancedSceneManager.Core.Runtime.isBuildMode","nameWithType":"Runtime.isBuildMode"},{"uid":"AdvancedSceneManager.Core.Runtime.wasStartedAsBuild","name":"wasStartedAsBuild","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_wasStartedAsBuild","commentId":"P:AdvancedSceneManager.Core.Runtime.wasStartedAsBuild","fullName":"AdvancedSceneManager.Core.Runtime.wasStartedAsBuild","nameWithType":"Runtime.wasStartedAsBuild"},{"uid":"AdvancedSceneManager.Core.Runtime.Start(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean)","name":"Start(SceneCollection, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Start_AdvancedSceneManager_Models_SceneCollection_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Runtime.Start(AdvancedSceneManager.Models.SceneCollection,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Core.Runtime.Start(AdvancedSceneManager.Models.SceneCollection, System.Boolean, System.Boolean)","nameWithType":"Runtime.Start(SceneCollection, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Core.Runtime.Restart(System.Boolean)","name":"Restart(Boolean)","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Restart_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.Runtime.Restart(System.Boolean)","fullName":"AdvancedSceneManager.Core.Runtime.Restart(System.Boolean)","nameWithType":"Runtime.Restart(Boolean)"},{"uid":"AdvancedSceneManager.Core.Runtime.RegisterQuitCallback(System.Collections.IEnumerator)","name":"RegisterQuitCallback(IEnumerator)","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_RegisterQuitCallback_System_Collections_IEnumerator_","commentId":"M:AdvancedSceneManager.Core.Runtime.RegisterQuitCallback(System.Collections.IEnumerator)","fullName":"AdvancedSceneManager.Core.Runtime.RegisterQuitCallback(System.Collections.IEnumerator)","nameWithType":"Runtime.RegisterQuitCallback(IEnumerator)"},{"uid":"AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback(System.Collections.IEnumerator)","name":"UnregisterQuitCallback(IEnumerator)","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_UnregisterQuitCallback_System_Collections_IEnumerator_","commentId":"M:AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback(System.Collections.IEnumerator)","fullName":"AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback(System.Collections.IEnumerator)","nameWithType":"Runtime.UnregisterQuitCallback(IEnumerator)"},{"uid":"AdvancedSceneManager.Core.Runtime.CancelQuit","name":"CancelQuit()","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_CancelQuit","commentId":"M:AdvancedSceneManager.Core.Runtime.CancelQuit","fullName":"AdvancedSceneManager.Core.Runtime.CancelQuit()","nameWithType":"Runtime.CancelQuit()"},{"uid":"AdvancedSceneManager.Core.Runtime.isQuitting","name":"isQuitting","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isQuitting","commentId":"P:AdvancedSceneManager.Core.Runtime.isQuitting","fullName":"AdvancedSceneManager.Core.Runtime.isQuitting","nameWithType":"Runtime.isQuitting"},{"uid":"AdvancedSceneManager.Core.Runtime.Quit(System.Boolean,System.Nullable{UnityEngine.Color},System.Single)","name":"Quit(Boolean, Nullable<Color>, Single)","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Quit_System_Boolean_System_Nullable_UnityEngine_Color__System_Single_","commentId":"M:AdvancedSceneManager.Core.Runtime.Quit(System.Boolean,System.Nullable{UnityEngine.Color},System.Single)","name.vb":"Quit(Boolean, Nullable(Of Color), Single)","fullName":"AdvancedSceneManager.Core.Runtime.Quit(System.Boolean, System.Nullable<UnityEngine.Color>, System.Single)","fullName.vb":"AdvancedSceneManager.Core.Runtime.Quit(System.Boolean, System.Nullable(Of UnityEngine.Color), System.Single)","nameWithType":"Runtime.Quit(Boolean, Nullable<Color>, Single)","nameWithType.vb":"Runtime.Quit(Boolean, Nullable(Of Color), Single)"},{"uid":"AdvancedSceneManager.Core.Runtime.isInitialized*","name":"isInitialized","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isInitialized_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.isInitialized","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.isInitialized","nameWithType":"Runtime.isInitialized"},{"uid":"AdvancedSceneManager.Core.Runtime.isBuildMode*","name":"isBuildMode","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isBuildMode_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.isBuildMode","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.isBuildMode","nameWithType":"Runtime.isBuildMode"},{"uid":"AdvancedSceneManager.Core.Runtime.wasStartedAsBuild*","name":"wasStartedAsBuild","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_wasStartedAsBuild_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.wasStartedAsBuild","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.wasStartedAsBuild","nameWithType":"Runtime.wasStartedAsBuild"},{"uid":"AdvancedSceneManager.Core.Runtime.Start*","name":"Start","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Start_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.Start","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.Start","nameWithType":"Runtime.Start"},{"uid":"AdvancedSceneManager.Core.Runtime.Restart*","name":"Restart","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Restart_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.Restart","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.Restart","nameWithType":"Runtime.Restart"},{"uid":"AdvancedSceneManager.Core.Runtime.RegisterQuitCallback*","name":"RegisterQuitCallback","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_RegisterQuitCallback_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.RegisterQuitCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.RegisterQuitCallback","nameWithType":"Runtime.RegisterQuitCallback"},{"uid":"AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback*","name":"UnregisterQuitCallback","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_UnregisterQuitCallback_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.UnregisterQuitCallback","nameWithType":"Runtime.UnregisterQuitCallback"},{"uid":"AdvancedSceneManager.Core.Runtime.CancelQuit*","name":"CancelQuit","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_CancelQuit_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.CancelQuit","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.CancelQuit","nameWithType":"Runtime.CancelQuit"},{"uid":"AdvancedSceneManager.Core.Runtime.isQuitting*","name":"isQuitting","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_isQuitting_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.isQuitting","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.isQuitting","nameWithType":"Runtime.isQuitting"},{"uid":"AdvancedSceneManager.Core.Runtime.Quit*","name":"Quit","href":"~/api/AdvancedSceneManager.Core.Runtime.yml#AdvancedSceneManager_Core_Runtime_Quit_","commentId":"Overload:AdvancedSceneManager.Core.Runtime.Quit","isSpec":"True","fullName":"AdvancedSceneManager.Core.Runtime.Quit","nameWithType":"Runtime.Quit"}],"api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen","name":"PressAnyButtonLoadingScreen","href":"~/api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen","fullName":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen","nameWithType":"PressAnyButtonLoadingScreen"},{"uid":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml#AdvancedSceneManager_Defaults_PressAnyButtonLoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"PressAnyButtonLoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml#AdvancedSceneManager_Defaults_PressAnyButtonLoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"PressAnyButtonLoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml#AdvancedSceneManager_Defaults_PressAnyButtonLoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnOpen","nameWithType":"PressAnyButtonLoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.yml#AdvancedSceneManager_Defaults_PressAnyButtonLoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.PressAnyButtonLoadingScreen.OnClose","nameWithType":"PressAnyButtonLoadingScreen.OnClose"}],"api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen","name":"QuoteLoadingScreen","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.QuoteLoadingScreen","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen","nameWithType":"QuoteLoadingScreen"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.quotes","name":"quotes","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_quotes","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.quotes","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.quotes","nameWithType":"QuoteLoadingScreen.quotes"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Background","name":"Background","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_Background","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.Background","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Background","nameWithType":"QuoteLoadingScreen.Background"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.fade","name":"fade","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_fade","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.fade","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.fade","nameWithType":"QuoteLoadingScreen.fade"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Quote","name":"Quote","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_Quote","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.Quote","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Quote","nameWithType":"QuoteLoadingScreen.Quote"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Name","name":"Name","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_Name","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.Name","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.Name","nameWithType":"QuoteLoadingScreen.Name"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.fadeDuration","name":"fadeDuration","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_fadeDuration","commentId":"F:AdvancedSceneManager.Defaults.QuoteLoadingScreen.fadeDuration","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.fadeDuration","nameWithType":"QuoteLoadingScreen.fadeDuration"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"QuoteLoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"QuoteLoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnOpen","nameWithType":"QuoteLoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Defaults.QuoteLoadingScreen.yml#AdvancedSceneManager_Defaults_QuoteLoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.QuoteLoadingScreen.OnClose","nameWithType":"QuoteLoadingScreen.OnClose"}],"api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml":[{"uid":"AdvancedSceneManager.Editor.IUIToolkitEditor","name":"IUIToolkitEditor","href":"~/api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml","commentId":"T:AdvancedSceneManager.Editor.IUIToolkitEditor","fullName":"AdvancedSceneManager.Editor.IUIToolkitEditor","nameWithType":"IUIToolkitEditor"},{"uid":"AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml#AdvancedSceneManager_Editor_IUIToolkitEditor_rootVisualElement","commentId":"P:AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement","fullName":"AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement","nameWithType":"IUIToolkitEditor.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.IUIToolkitEditor.position","name":"position","href":"~/api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml#AdvancedSceneManager_Editor_IUIToolkitEditor_position","commentId":"P:AdvancedSceneManager.Editor.IUIToolkitEditor.position","fullName":"AdvancedSceneManager.Editor.IUIToolkitEditor.position","nameWithType":"IUIToolkitEditor.position"},{"uid":"AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement*","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml#AdvancedSceneManager_Editor_IUIToolkitEditor_rootVisualElement_","commentId":"Overload:AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement","isSpec":"True","fullName":"AdvancedSceneManager.Editor.IUIToolkitEditor.rootVisualElement","nameWithType":"IUIToolkitEditor.rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.IUIToolkitEditor.position*","name":"position","href":"~/api/AdvancedSceneManager.Editor.IUIToolkitEditor.yml#AdvancedSceneManager_Editor_IUIToolkitEditor_position_","commentId":"Overload:AdvancedSceneManager.Editor.IUIToolkitEditor.position","isSpec":"True","fullName":"AdvancedSceneManager.Editor.IUIToolkitEditor.position","nameWithType":"IUIToolkitEditor.position"}],"api/AdvancedSceneManager.Editor.ObjectField.UxmlFactory.yml":[{"uid":"AdvancedSceneManager.Editor.ObjectField.UxmlFactory","name":"ObjectField.UxmlFactory","href":"~/api/AdvancedSceneManager.Editor.ObjectField.UxmlFactory.yml","commentId":"T:AdvancedSceneManager.Editor.ObjectField.UxmlFactory","fullName":"AdvancedSceneManager.Editor.ObjectField.UxmlFactory","nameWithType":"ObjectField.UxmlFactory"}],"api/AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.yml":[{"uid":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent","name":"SceneField.SceneChangedEvent","href":"~/api/AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.yml","commentId":"T:AdvancedSceneManager.Editor.SceneField.SceneChangedEvent","fullName":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent","nameWithType":"SceneField.SceneChangedEvent"},{"uid":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.Scene)","name":"SceneChangedEvent(Scene, Scene)","href":"~/api/AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.yml#AdvancedSceneManager_Editor_SceneField_SceneChangedEvent__ctor_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.SceneChangedEvent(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.Scene)","nameWithType":"SceneField.SceneChangedEvent.SceneChangedEvent(Scene, Scene)"},{"uid":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.#ctor*","name":"SceneChangedEvent","href":"~/api/AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.yml#AdvancedSceneManager_Editor_SceneField_SceneChangedEvent__ctor_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.SceneChangedEvent.SceneChangedEvent","nameWithType":"SceneField.SceneChangedEvent.SceneChangedEvent"}],"api/AdvancedSceneManager.Editor.SceneField.UxmlFactory.yml":[{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlFactory","name":"SceneField.UxmlFactory","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlFactory.yml","commentId":"T:AdvancedSceneManager.Editor.SceneField.UxmlFactory","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlFactory","nameWithType":"SceneField.UxmlFactory"}],"api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml":[{"uid":"AdvancedSceneManager.Editor.ScenePropertyDrawer","name":"ScenePropertyDrawer","href":"~/api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml","commentId":"T:AdvancedSceneManager.Editor.ScenePropertyDrawer","fullName":"AdvancedSceneManager.Editor.ScenePropertyDrawer","nameWithType":"ScenePropertyDrawer"},{"uid":"AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI(UnityEngine.Rect,UnityEditor.SerializedProperty,UnityEngine.GUIContent)","name":"OnGUI(Rect, SerializedProperty, GUIContent)","href":"~/api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml#AdvancedSceneManager_Editor_ScenePropertyDrawer_OnGUI_UnityEngine_Rect_UnityEditor_SerializedProperty_UnityEngine_GUIContent_","commentId":"M:AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI(UnityEngine.Rect,UnityEditor.SerializedProperty,UnityEngine.GUIContent)","fullName":"AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI(UnityEngine.Rect, UnityEditor.SerializedProperty, UnityEngine.GUIContent)","nameWithType":"ScenePropertyDrawer.OnGUI(Rect, SerializedProperty, GUIContent)"},{"uid":"AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField``1(UnityEngine.Rect,``0,System.Func{UnityEngine.Object,System.ValueTuple{``0,System.Boolean}},System.Type[])","name":"ObjectField<T>(Rect, T, Func<Object, (T obj, Boolean didConvert)>, Type[])","href":"~/api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml#AdvancedSceneManager_Editor_ScenePropertyDrawer_ObjectField__1_UnityEngine_Rect___0_System_Func_UnityEngine_Object_System_ValueTuple___0_System_Boolean___System_Type___","commentId":"M:AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField``1(UnityEngine.Rect,``0,System.Func{UnityEngine.Object,System.ValueTuple{``0,System.Boolean}},System.Type[])","name.vb":"ObjectField(Of T)(Rect, T, Func(Of Object, (obj As T, didConvert As Boolean)(Of T, Boolean)), Type())","fullName":"AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField<T>(UnityEngine.Rect, T, System.Func<UnityEngine.Object, System.ValueTuple<T, System.Boolean>>, System.Type[])","fullName.vb":"AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField(Of T)(UnityEngine.Rect, T, System.Func(Of UnityEngine.Object, System.ValueTuple(Of T, System.Boolean)), System.Type())","nameWithType":"ScenePropertyDrawer.ObjectField<T>(Rect, T, Func<Object, (T obj, Boolean didConvert)>, Type[])","nameWithType.vb":"ScenePropertyDrawer.ObjectField(Of T)(Rect, T, Func(Of Object, (obj As T, didConvert As Boolean)(Of T, Boolean)), Type())"},{"uid":"AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI*","name":"OnGUI","href":"~/api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml#AdvancedSceneManager_Editor_ScenePropertyDrawer_OnGUI_","commentId":"Overload:AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenePropertyDrawer.OnGUI","nameWithType":"ScenePropertyDrawer.OnGUI"},{"uid":"AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField*","name":"ObjectField","href":"~/api/AdvancedSceneManager.Editor.ScenePropertyDrawer.yml#AdvancedSceneManager_Editor_ScenePropertyDrawer_ObjectField_","commentId":"Overload:AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenePropertyDrawer.ObjectField","nameWithType":"ScenePropertyDrawer.ObjectField"}],"api/AdvancedSceneManager.Editor.ScenesTab.yml":[{"uid":"AdvancedSceneManager.Editor.ScenesTab","name":"ScenesTab","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml","commentId":"T:AdvancedSceneManager.Editor.ScenesTab","fullName":"AdvancedSceneManager.Editor.ScenesTab","nameWithType":"ScenesTab"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnEnable(UnityEngine.UIElements.VisualElement)","name":"OnEnable(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnEnable_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.OnEnable(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnEnable(UnityEngine.UIElements.VisualElement)","nameWithType":"ScenesTab.OnEnable(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnDisable","name":"OnDisable()","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnDisable","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.OnDisable","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnDisable()","nameWithType":"ScenesTab.OnDisable()"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.Open(System.ValueTuple{AdvancedSceneManager.Models.SceneCollection,System.Int32},System.Boolean)","name":"Open((SceneCollection collection, Int32 i), Boolean)","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_Open_System_ValueTuple_AdvancedSceneManager_Models_SceneCollection_System_Int32__System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.Open(System.ValueTuple{AdvancedSceneManager.Models.SceneCollection,System.Int32},System.Boolean)","name.vb":"Open((collection As SceneCollection, i As Int32)(Of SceneCollection, Int32), Boolean)","fullName":"AdvancedSceneManager.Editor.ScenesTab.Open(System.ValueTuple<AdvancedSceneManager.Models.SceneCollection, System.Int32>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.ScenesTab.Open(System.ValueTuple(Of AdvancedSceneManager.Models.SceneCollection, System.Int32), System.Boolean)","nameWithType":"ScenesTab.Open((SceneCollection collection, Int32 i), Boolean)","nameWithType.vb":"ScenesTab.Open((collection As SceneCollection, i As Int32)(Of SceneCollection, Int32), Boolean)"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.Path(System.ValueTuple{AdvancedSceneManager.Models.SceneCollection,System.Int32})","name":"Path((SceneCollection collection, Int32 i))","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_Path_System_ValueTuple_AdvancedSceneManager_Models_SceneCollection_System_Int32__","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.Path(System.ValueTuple{AdvancedSceneManager.Models.SceneCollection,System.Int32})","name.vb":"Path((collection As SceneCollection, i As Int32)(Of SceneCollection, Int32))","fullName":"AdvancedSceneManager.Editor.ScenesTab.Path(System.ValueTuple<AdvancedSceneManager.Models.SceneCollection, System.Int32>)","fullName.vb":"AdvancedSceneManager.Editor.ScenesTab.Path(System.ValueTuple(Of AdvancedSceneManager.Models.SceneCollection, System.Int32))","nameWithType":"ScenesTab.Path((SceneCollection collection, Int32 i))","nameWithType.vb":"ScenesTab.Path((collection As SceneCollection, i As Int32)(Of SceneCollection, Int32))"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.FooterButtons","name":"FooterButtons","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_FooterButtons","commentId":"P:AdvancedSceneManager.Editor.ScenesTab.FooterButtons","fullName":"AdvancedSceneManager.Editor.ScenesTab.FooterButtons","nameWithType":"ScenesTab.FooterButtons"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnReorderStart(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement)","name":"OnReorderStart(SceneManagerWindow.DragAndDropReorder.DragElement)","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnReorderStart_AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.OnReorderStart(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement)","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnReorderStart(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement)","nameWithType":"ScenesTab.OnReorderStart(SceneManagerWindow.DragAndDropReorder.DragElement)"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement,System.Int32)","name":"OnReorderEnd(SceneManagerWindow.DragAndDropReorder.DragElement, Int32)","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnReorderEnd_AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement,System.Int32)","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement, System.Int32)","nameWithType":"ScenesTab.OnReorderEnd(SceneManagerWindow.DragAndDropReorder.DragElement, Int32)"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnEnable","nameWithType":"ScenesTab.OnEnable"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnDisable*","name":"OnDisable","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnDisable_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.OnDisable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnDisable","nameWithType":"ScenesTab.OnDisable"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_Open_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.Open","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.Open","nameWithType":"ScenesTab.Open"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.Path*","name":"Path","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_Path_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.Path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.Path","nameWithType":"ScenesTab.Path"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.FooterButtons*","name":"FooterButtons","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_FooterButtons_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.FooterButtons","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.FooterButtons","nameWithType":"ScenesTab.FooterButtons"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnReorderStart*","name":"OnReorderStart","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnReorderStart_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.OnReorderStart","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnReorderStart","nameWithType":"ScenesTab.OnReorderStart"},{"uid":"AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd*","name":"OnReorderEnd","href":"~/api/AdvancedSceneManager.Editor.ScenesTab.yml#AdvancedSceneManager_Editor_ScenesTab_OnReorderEnd_","commentId":"Overload:AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd","isSpec":"True","fullName":"AdvancedSceneManager.Editor.ScenesTab.OnReorderEnd","nameWithType":"ScenesTab.OnReorderEnd"}],"api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt","name":"EditorGUIUtilityExt","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt","fullName":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt","nameWithType":"EditorGUIUtilityExt"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset(UnityEngine.Object,System.Int32)","name":"PingOrOpenAsset(Object, Int32)","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml#AdvancedSceneManager_Editor_Utility_EditorGUIUtilityExt_PingOrOpenAsset_UnityEngine_Object_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset(UnityEngine.Object,System.Int32)","fullName":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset(UnityEngine.Object, System.Int32)","nameWithType":"EditorGUIUtilityExt.PingOrOpenAsset(Object, Int32)"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor","name":"GetDefaultBackgroundColor()","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml#AdvancedSceneManager_Editor_Utility_EditorGUIUtilityExt_GetDefaultBackgroundColor","commentId":"M:AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor","fullName":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor()","nameWithType":"EditorGUIUtilityExt.GetDefaultBackgroundColor()"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset*","name":"PingOrOpenAsset","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml#AdvancedSceneManager_Editor_Utility_EditorGUIUtilityExt_PingOrOpenAsset_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.PingOrOpenAsset","nameWithType":"EditorGUIUtilityExt.PingOrOpenAsset"},{"uid":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor*","name":"GetDefaultBackgroundColor","href":"~/api/AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.yml#AdvancedSceneManager_Editor_Utility_EditorGUIUtilityExt_GetDefaultBackgroundColor_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.EditorGUIUtilityExt.GetDefaultBackgroundColor","nameWithType":"EditorGUIUtilityExt.GetDefaultBackgroundColor"}],"api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2","name":"GenericPrompt<T, TSelf>","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.GenericPrompt`2","name.vb":"GenericPrompt(Of T, TSelf)","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf)","nameWithType":"GenericPrompt<T, TSelf>","nameWithType.vb":"GenericPrompt(Of T, TSelf)"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.validate","name":"validate","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_validate","commentId":"F:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.validate","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.validate","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).validate","nameWithType":"GenericPrompt<T, TSelf>.validate","nameWithType.vb":"GenericPrompt(Of T, TSelf).validate"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Validate(`0)","name":"Validate(T)","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_Validate__0_","commentId":"M:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Validate(`0)","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.Validate(T)","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).Validate(T)","nameWithType":"GenericPrompt<T, TSelf>.Validate(T)","nameWithType.vb":"GenericPrompt(Of T, TSelf).Validate(T)"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Prompt(`0,System.Func{`0,System.ValueTuple{System.Boolean,System.String}}[])","name":"Prompt(T, Func<T, (Boolean isValid, String message)>[])","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_Prompt__0_System_Func__0_System_ValueTuple_System_Boolean_System_String_____","commentId":"M:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Prompt(`0,System.Func{`0,System.ValueTuple{System.Boolean,System.String}}[])","name.vb":"Prompt(T, Func(Of T, (isValid As Boolean, message As String)(Of Boolean, String))())","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.Prompt(T, System.Func<T, System.ValueTuple<System.Boolean, System.String>>[])","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).Prompt(T, System.Func(Of T, System.ValueTuple(Of System.Boolean, System.String))())","nameWithType":"GenericPrompt<T, TSelf>.Prompt(T, Func<T, (Boolean isValid, String message)>[])","nameWithType.vb":"GenericPrompt(Of T, TSelf).Prompt(T, Func(Of T, (isValid As Boolean, message As String)(Of Boolean, String))())"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.OnContentGUI(`0@)","name":"OnContentGUI(ref T)","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_OnContentGUI__0__","commentId":"M:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.OnContentGUI(`0@)","name.vb":"OnContentGUI(ByRef T)","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.OnContentGUI(ref T)","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).OnContentGUI(ByRef T)","nameWithType":"GenericPrompt<T, TSelf>.OnContentGUI(ref T)","nameWithType.vb":"GenericPrompt(Of T, TSelf).OnContentGUI(ByRef T)"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_title","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.title","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.title","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).title","nameWithType":"GenericPrompt<T, TSelf>.title","nameWithType.vb":"GenericPrompt(Of T, TSelf).title"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.updateSizeAutomatically","name":"updateSizeAutomatically","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_updateSizeAutomatically","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.updateSizeAutomatically","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.updateSizeAutomatically","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).updateSizeAutomatically","nameWithType":"GenericPrompt<T, TSelf>.updateSizeAutomatically","nameWithType.vb":"GenericPrompt(Of T, TSelf).updateSizeAutomatically"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.extraHeight","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_extraHeight","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.extraHeight","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.extraHeight","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).extraHeight","nameWithType":"GenericPrompt<T, TSelf>.extraHeight","nameWithType.vb":"GenericPrompt(Of T, TSelf).extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.width","name":"width","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_width","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.width","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.width","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).width","nameWithType":"GenericPrompt<T, TSelf>.width","nameWithType.vb":"GenericPrompt(Of T, TSelf).width"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.okButton","name":"okButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_okButton","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.okButton","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.okButton","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).okButton","nameWithType":"GenericPrompt<T, TSelf>.okButton","nameWithType.vb":"GenericPrompt(Of T, TSelf).okButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.cancelButton","name":"cancelButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_cancelButton","commentId":"P:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.cancelButton","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.cancelButton","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).cancelButton","nameWithType":"GenericPrompt<T, TSelf>.cancelButton","nameWithType.vb":"GenericPrompt(Of T, TSelf).cancelButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Validate*","name":"Validate","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_Validate_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Validate","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.Validate","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).Validate","nameWithType":"GenericPrompt<T, TSelf>.Validate","nameWithType.vb":"GenericPrompt(Of T, TSelf).Validate"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Prompt*","name":"Prompt","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_Prompt_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.Prompt","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.Prompt","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).Prompt","nameWithType":"GenericPrompt<T, TSelf>.Prompt","nameWithType.vb":"GenericPrompt(Of T, TSelf).Prompt"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.OnContentGUI","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).OnContentGUI","nameWithType":"GenericPrompt<T, TSelf>.OnContentGUI","nameWithType.vb":"GenericPrompt(Of T, TSelf).OnContentGUI"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.title","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).title","nameWithType":"GenericPrompt<T, TSelf>.title","nameWithType.vb":"GenericPrompt(Of T, TSelf).title"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.updateSizeAutomatically*","name":"updateSizeAutomatically","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_updateSizeAutomatically_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.updateSizeAutomatically","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.updateSizeAutomatically","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).updateSizeAutomatically","nameWithType":"GenericPrompt<T, TSelf>.updateSizeAutomatically","nameWithType.vb":"GenericPrompt(Of T, TSelf).updateSizeAutomatically"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.extraHeight*","name":"extraHeight","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_extraHeight_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.extraHeight","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.extraHeight","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).extraHeight","nameWithType":"GenericPrompt<T, TSelf>.extraHeight","nameWithType.vb":"GenericPrompt(Of T, TSelf).extraHeight"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.width*","name":"width","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_width_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.width","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.width","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).width","nameWithType":"GenericPrompt<T, TSelf>.width","nameWithType.vb":"GenericPrompt(Of T, TSelf).width"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.okButton*","name":"okButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_okButton_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.okButton","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.okButton","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).okButton","nameWithType":"GenericPrompt<T, TSelf>.okButton","nameWithType.vb":"GenericPrompt(Of T, TSelf).okButton"},{"uid":"AdvancedSceneManager.Editor.Utility.GenericPrompt`2.cancelButton*","name":"cancelButton","href":"~/api/AdvancedSceneManager.Editor.Utility.GenericPrompt-2.yml#AdvancedSceneManager_Editor_Utility_GenericPrompt_2_cancelButton_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.GenericPrompt`2.cancelButton","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.GenericPrompt<T, TSelf>.cancelButton","fullName.vb":"AdvancedSceneManager.Editor.Utility.GenericPrompt(Of T, TSelf).cancelButton","nameWithType":"GenericPrompt<T, TSelf>.cancelButton","nameWithType.vb":"GenericPrompt(Of T, TSelf).cancelButton"}],"api/AdvancedSceneManager.Editor.Utility.PromptInt.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt","name":"PromptInt","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PromptInt","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt","nameWithType":"PromptInt"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_title","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptInt.title","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.title","nameWithType":"PromptInt.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.Validate(System.String)","name":"Validate(String)","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_Validate_System_String_","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptInt.Validate(System.String)","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.Validate(System.String)","nameWithType":"PromptInt.Validate(String)"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI(System.String@)","name":"OnContentGUI(ref String)","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_OnContentGUI_System_String__","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI(System.String@)","name.vb":"OnContentGUI(ByRef String)","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI(ref System.String)","fullName.vb":"AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI(ByRef System.String)","nameWithType":"PromptInt.OnContentGUI(ref String)","nameWithType.vb":"PromptInt.OnContentGUI(ByRef String)"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptInt.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.title","nameWithType":"PromptInt.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.Validate*","name":"Validate","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_Validate_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptInt.Validate","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.Validate","nameWithType":"PromptInt.Validate"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptInt.yml#AdvancedSceneManager_Editor_Utility_PromptInt_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptInt.OnContentGUI","nameWithType":"PromptInt.OnContentGUI"}],"api/AdvancedSceneManager.Editor.Utility.PromptKey.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.PromptKey","name":"PromptKey","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptKey.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.PromptKey","fullName":"AdvancedSceneManager.Editor.Utility.PromptKey","nameWithType":"PromptKey"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptKey.title","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptKey.yml#AdvancedSceneManager_Editor_Utility_PromptKey_title","commentId":"P:AdvancedSceneManager.Editor.Utility.PromptKey.title","fullName":"AdvancedSceneManager.Editor.Utility.PromptKey.title","nameWithType":"PromptKey.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI(System.ValueTuple{UnityEngine.EventModifiers,UnityEngine.KeyCode}@)","name":"OnContentGUI(ref (EventModifiers modifiers, KeyCode key))","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptKey.yml#AdvancedSceneManager_Editor_Utility_PromptKey_OnContentGUI_System_ValueTuple_UnityEngine_EventModifiers_UnityEngine_KeyCode___","commentId":"M:AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI(System.ValueTuple{UnityEngine.EventModifiers,UnityEngine.KeyCode}@)","name.vb":"OnContentGUI(ByRef (modifiers As EventModifiers, key As KeyCode)(Of EventModifiers, KeyCode))","fullName":"AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI(ref System.ValueTuple<UnityEngine.EventModifiers, UnityEngine.KeyCode>)","fullName.vb":"AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI(ByRef System.ValueTuple(Of UnityEngine.EventModifiers, UnityEngine.KeyCode))","nameWithType":"PromptKey.OnContentGUI(ref (EventModifiers modifiers, KeyCode key))","nameWithType.vb":"PromptKey.OnContentGUI(ByRef (modifiers As EventModifiers, key As KeyCode)(Of EventModifiers, KeyCode))"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptKey.title*","name":"title","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptKey.yml#AdvancedSceneManager_Editor_Utility_PromptKey_title_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptKey.title","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptKey.title","nameWithType":"PromptKey.title"},{"uid":"AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI*","name":"OnContentGUI","href":"~/api/AdvancedSceneManager.Editor.Utility.PromptKey.yml#AdvancedSceneManager_Editor_Utility_PromptKey_OnContentGUI_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.PromptKey.OnContentGUI","nameWithType":"PromptKey.OnContentGUI"}],"api/AdvancedSceneManager.Exceptions.OpenSceneException.yml":[{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException","name":"OpenSceneException","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml","commentId":"T:AdvancedSceneManager.Exceptions.OpenSceneException","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException","nameWithType":"OpenSceneException"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection,System.String)","name":"OpenSceneException(Scene, SceneCollection, String)","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException__ctor_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneCollection_System_String_","commentId":"M:AdvancedSceneManager.Exceptions.OpenSceneException.#ctor(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneCollection,System.String)","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.OpenSceneException(AdvancedSceneManager.Models.Scene, AdvancedSceneManager.Models.SceneCollection, System.String)","nameWithType":"OpenSceneException.OpenSceneException(Scene, SceneCollection, String)"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.collection","name":"collection","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException_collection","commentId":"P:AdvancedSceneManager.Exceptions.OpenSceneException.collection","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.collection","nameWithType":"OpenSceneException.collection"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.scene","name":"scene","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException_scene","commentId":"P:AdvancedSceneManager.Exceptions.OpenSceneException.scene","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.scene","nameWithType":"OpenSceneException.scene"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.#ctor*","name":"OpenSceneException","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException__ctor_","commentId":"Overload:AdvancedSceneManager.Exceptions.OpenSceneException.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.OpenSceneException","nameWithType":"OpenSceneException.OpenSceneException"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.collection*","name":"collection","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException_collection_","commentId":"Overload:AdvancedSceneManager.Exceptions.OpenSceneException.collection","isSpec":"True","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.collection","nameWithType":"OpenSceneException.collection"},{"uid":"AdvancedSceneManager.Exceptions.OpenSceneException.scene*","name":"scene","href":"~/api/AdvancedSceneManager.Exceptions.OpenSceneException.yml#AdvancedSceneManager_Exceptions_OpenSceneException_scene_","commentId":"Overload:AdvancedSceneManager.Exceptions.OpenSceneException.scene","isSpec":"True","fullName":"AdvancedSceneManager.Exceptions.OpenSceneException.scene","nameWithType":"OpenSceneException.scene"}],"api/AdvancedSceneManager.Exceptions.yml":[{"uid":"AdvancedSceneManager.Exceptions","name":"AdvancedSceneManager.Exceptions","href":"~/api/AdvancedSceneManager.Exceptions.yml","commentId":"N:AdvancedSceneManager.Exceptions","fullName":"AdvancedSceneManager.Exceptions","nameWithType":"AdvancedSceneManager.Exceptions"}],"api/AdvancedSceneManager.Models.IsOpenReturnValue.yml":[{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue","name":"IsOpenReturnValue","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml","commentId":"T:AdvancedSceneManager.Models.IsOpenReturnValue","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue","nameWithType":"IsOpenReturnValue"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.withCollection","name":"withCollection","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_withCollection","commentId":"F:AdvancedSceneManager.Models.IsOpenReturnValue.withCollection","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.withCollection","nameWithType":"IsOpenReturnValue.withCollection"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.asStandalone","name":"asStandalone","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_asStandalone","commentId":"F:AdvancedSceneManager.Models.IsOpenReturnValue.asStandalone","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.asStandalone","nameWithType":"IsOpenReturnValue.asStandalone"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.isPreloaded","name":"isPreloaded","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_isPreloaded","commentId":"F:AdvancedSceneManager.Models.IsOpenReturnValue.isPreloaded","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.isPreloaded","nameWithType":"IsOpenReturnValue.isPreloaded"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(AdvancedSceneManager.Models.IsOpenReturnValue)~System.Boolean","name":"Implicit(IsOpenReturnValue to Boolean)","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_op_Implicit_AdvancedSceneManager_Models_IsOpenReturnValue__System_Boolean","commentId":"M:AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(AdvancedSceneManager.Models.IsOpenReturnValue)~System.Boolean","name.vb":"Widening(IsOpenReturnValue to Boolean)","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.Implicit(AdvancedSceneManager.Models.IsOpenReturnValue to System.Boolean)","fullName.vb":"AdvancedSceneManager.Models.IsOpenReturnValue.Widening(AdvancedSceneManager.Models.IsOpenReturnValue to System.Boolean)","nameWithType":"IsOpenReturnValue.Implicit(IsOpenReturnValue to Boolean)","nameWithType.vb":"IsOpenReturnValue.Widening(IsOpenReturnValue to Boolean)"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(System.ValueTuple{System.Boolean,System.Boolean})~AdvancedSceneManager.Models.IsOpenReturnValue","name":"Implicit((Boolean withCollection, Boolean asStandalone) to IsOpenReturnValue)","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_op_Implicit_System_ValueTuple_System_Boolean_System_Boolean___AdvancedSceneManager_Models_IsOpenReturnValue","commentId":"M:AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(System.ValueTuple{System.Boolean,System.Boolean})~AdvancedSceneManager.Models.IsOpenReturnValue","name.vb":"Widening((withCollection As Boolean, asStandalone As Boolean)(Of Boolean, Boolean) to IsOpenReturnValue)","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.Implicit(System.ValueTuple<System.Boolean, System.Boolean> to AdvancedSceneManager.Models.IsOpenReturnValue)","fullName.vb":"AdvancedSceneManager.Models.IsOpenReturnValue.Widening(System.ValueTuple(Of System.Boolean, System.Boolean) to AdvancedSceneManager.Models.IsOpenReturnValue)","nameWithType":"IsOpenReturnValue.Implicit((Boolean withCollection, Boolean asStandalone) to IsOpenReturnValue)","nameWithType.vb":"IsOpenReturnValue.Widening((withCollection As Boolean, asStandalone As Boolean)(Of Boolean, Boolean) to IsOpenReturnValue)"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(System.ValueTuple{System.Boolean,System.Boolean,System.Boolean})~AdvancedSceneManager.Models.IsOpenReturnValue","name":"Implicit((Boolean withCollection, Boolean asStandalone, Boolean isPreloaded) to IsOpenReturnValue)","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_op_Implicit_System_ValueTuple_System_Boolean_System_Boolean_System_Boolean___AdvancedSceneManager_Models_IsOpenReturnValue","commentId":"M:AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit(System.ValueTuple{System.Boolean,System.Boolean,System.Boolean})~AdvancedSceneManager.Models.IsOpenReturnValue","name.vb":"Widening((withCollection As Boolean, asStandalone As Boolean, isPreloaded As Boolean)(Of Boolean, Boolean, Boolean) to IsOpenReturnValue)","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.Implicit(System.ValueTuple<System.Boolean, System.Boolean, System.Boolean> to AdvancedSceneManager.Models.IsOpenReturnValue)","fullName.vb":"AdvancedSceneManager.Models.IsOpenReturnValue.Widening(System.ValueTuple(Of System.Boolean, System.Boolean, System.Boolean) to AdvancedSceneManager.Models.IsOpenReturnValue)","nameWithType":"IsOpenReturnValue.Implicit((Boolean withCollection, Boolean asStandalone, Boolean isPreloaded) to IsOpenReturnValue)","nameWithType.vb":"IsOpenReturnValue.Widening((withCollection As Boolean, asStandalone As Boolean, isPreloaded As Boolean)(Of Boolean, Boolean, Boolean) to IsOpenReturnValue)"},{"uid":"AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit*","name":"Implicit","href":"~/api/AdvancedSceneManager.Models.IsOpenReturnValue.yml#AdvancedSceneManager_Models_IsOpenReturnValue_op_Implicit_","commentId":"Overload:AdvancedSceneManager.Models.IsOpenReturnValue.op_Implicit","isSpec":"True","name.vb":"Widening","fullName":"AdvancedSceneManager.Models.IsOpenReturnValue.Implicit","fullName.vb":"AdvancedSceneManager.Models.IsOpenReturnValue.Widening","nameWithType":"IsOpenReturnValue.Implicit","nameWithType.vb":"IsOpenReturnValue.Widening"}],"api/AdvancedSceneManager.Models.LoadingScreenUsage.yml":[{"uid":"AdvancedSceneManager.Models.LoadingScreenUsage","name":"LoadingScreenUsage","href":"~/api/AdvancedSceneManager.Models.LoadingScreenUsage.yml","commentId":"T:AdvancedSceneManager.Models.LoadingScreenUsage","fullName":"AdvancedSceneManager.Models.LoadingScreenUsage","nameWithType":"LoadingScreenUsage"},{"uid":"AdvancedSceneManager.Models.LoadingScreenUsage.DoNotUse","name":"DoNotUse","href":"~/api/AdvancedSceneManager.Models.LoadingScreenUsage.yml#AdvancedSceneManager_Models_LoadingScreenUsage_DoNotUse","commentId":"F:AdvancedSceneManager.Models.LoadingScreenUsage.DoNotUse","fullName":"AdvancedSceneManager.Models.LoadingScreenUsage.DoNotUse","nameWithType":"LoadingScreenUsage.DoNotUse"},{"uid":"AdvancedSceneManager.Models.LoadingScreenUsage.UseDefault","name":"UseDefault","href":"~/api/AdvancedSceneManager.Models.LoadingScreenUsage.yml#AdvancedSceneManager_Models_LoadingScreenUsage_UseDefault","commentId":"F:AdvancedSceneManager.Models.LoadingScreenUsage.UseDefault","fullName":"AdvancedSceneManager.Models.LoadingScreenUsage.UseDefault","nameWithType":"LoadingScreenUsage.UseDefault"},{"uid":"AdvancedSceneManager.Models.LoadingScreenUsage.Override","name":"Override","href":"~/api/AdvancedSceneManager.Models.LoadingScreenUsage.yml#AdvancedSceneManager_Models_LoadingScreenUsage_Override","commentId":"F:AdvancedSceneManager.Models.LoadingScreenUsage.Override","fullName":"AdvancedSceneManager.Models.LoadingScreenUsage.Override","nameWithType":"LoadingScreenUsage.Override"}],"api/AdvancedSceneManager.Models.Profile.yml":[{"uid":"AdvancedSceneManager.Models.Profile","name":"Profile","href":"~/api/AdvancedSceneManager.Models.Profile.yml","commentId":"T:AdvancedSceneManager.Models.Profile","fullName":"AdvancedSceneManager.Models.Profile","nameWithType":"Profile"},{"uid":"AdvancedSceneManager.Models.Profile.FindAll","name":"FindAll()","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_FindAll","commentId":"M:AdvancedSceneManager.Models.Profile.FindAll","fullName":"AdvancedSceneManager.Models.Profile.FindAll()","nameWithType":"Profile.FindAll()"},{"uid":"AdvancedSceneManager.Models.Profile.Find(System.Func{AdvancedSceneManager.Models.Profile,System.Boolean})","name":"Find(Func<Profile, Boolean>)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Find_System_Func_AdvancedSceneManager_Models_Profile_System_Boolean__","commentId":"M:AdvancedSceneManager.Models.Profile.Find(System.Func{AdvancedSceneManager.Models.Profile,System.Boolean})","name.vb":"Find(Func(Of Profile, Boolean))","fullName":"AdvancedSceneManager.Models.Profile.Find(System.Func<AdvancedSceneManager.Models.Profile, System.Boolean>)","fullName.vb":"AdvancedSceneManager.Models.Profile.Find(System.Func(Of AdvancedSceneManager.Models.Profile, System.Boolean))","nameWithType":"Profile.Find(Func<Profile, Boolean>)","nameWithType.vb":"Profile.Find(Func(Of Profile, Boolean))"},{"uid":"AdvancedSceneManager.Models.Profile.Find(System.String)","name":"Find(String)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Find_System_String_","commentId":"M:AdvancedSceneManager.Models.Profile.Find(System.String)","fullName":"AdvancedSceneManager.Models.Profile.Find(System.String)","nameWithType":"Profile.Find(String)"},{"uid":"AdvancedSceneManager.Models.Profile.name","name":"name","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_name","commentId":"P:AdvancedSceneManager.Models.Profile.name","fullName":"AdvancedSceneManager.Models.Profile.name","nameWithType":"Profile.name"},{"uid":"AdvancedSceneManager.Models.Profile.MarkAsDirty","name":"MarkAsDirty()","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_MarkAsDirty","commentId":"M:AdvancedSceneManager.Models.Profile.MarkAsDirty","fullName":"AdvancedSceneManager.Models.Profile.MarkAsDirty()","nameWithType":"Profile.MarkAsDirty()"},{"uid":"AdvancedSceneManager.Models.Profile.current","name":"current","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_current","commentId":"P:AdvancedSceneManager.Models.Profile.current","fullName":"AdvancedSceneManager.Models.Profile.current","nameWithType":"Profile.current"},{"uid":"AdvancedSceneManager.Models.Profile.onProfileChanged","name":"onProfileChanged","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_onProfileChanged","commentId":"E:AdvancedSceneManager.Models.Profile.onProfileChanged","fullName":"AdvancedSceneManager.Models.Profile.onProfileChanged","nameWithType":"Profile.onProfileChanged"},{"uid":"AdvancedSceneManager.Models.Profile.collections","name":"collections","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_collections","commentId":"P:AdvancedSceneManager.Models.Profile.collections","fullName":"AdvancedSceneManager.Models.Profile.collections","nameWithType":"Profile.collections"},{"uid":"AdvancedSceneManager.Models.Profile.scenes","name":"scenes","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_scenes","commentId":"P:AdvancedSceneManager.Models.Profile.scenes","fullName":"AdvancedSceneManager.Models.Profile.scenes","nameWithType":"Profile.scenes"},{"uid":"AdvancedSceneManager.Models.Profile.scenePaths","name":"scenePaths","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_scenePaths","commentId":"P:AdvancedSceneManager.Models.Profile.scenePaths","fullName":"AdvancedSceneManager.Models.Profile.scenePaths","nameWithType":"Profile.scenePaths"},{"uid":"AdvancedSceneManager.Models.Profile.StartupCollections","name":"StartupCollections()","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_StartupCollections","commentId":"M:AdvancedSceneManager.Models.Profile.StartupCollections","fullName":"AdvancedSceneManager.Models.Profile.StartupCollections()","nameWithType":"Profile.StartupCollections()"},{"uid":"AdvancedSceneManager.Models.Profile.CreateCollection(System.String,System.Action{AdvancedSceneManager.Models.SceneCollection})","name":"CreateCollection(String, Action<SceneCollection>)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_CreateCollection_System_String_System_Action_AdvancedSceneManager_Models_SceneCollection__","commentId":"M:AdvancedSceneManager.Models.Profile.CreateCollection(System.String,System.Action{AdvancedSceneManager.Models.SceneCollection})","name.vb":"CreateCollection(String, Action(Of SceneCollection))","fullName":"AdvancedSceneManager.Models.Profile.CreateCollection(System.String, System.Action<AdvancedSceneManager.Models.SceneCollection>)","fullName.vb":"AdvancedSceneManager.Models.Profile.CreateCollection(System.String, System.Action(Of AdvancedSceneManager.Models.SceneCollection))","nameWithType":"Profile.CreateCollection(String, Action<SceneCollection>)","nameWithType.vb":"Profile.CreateCollection(String, Action(Of SceneCollection))"},{"uid":"AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.SceneCollection)","name":"Add(SceneCollection)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Add_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"Profile.Add(SceneCollection)"},{"uid":"AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.SceneCollection)","name":"Remove(SceneCollection)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Remove_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"Profile.Remove(SceneCollection)"},{"uid":"AdvancedSceneManager.Models.Profile.PropertyChanged","name":"PropertyChanged","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_PropertyChanged","commentId":"E:AdvancedSceneManager.Models.Profile.PropertyChanged","fullName":"AdvancedSceneManager.Models.Profile.PropertyChanged","nameWithType":"Profile.PropertyChanged"},{"uid":"AdvancedSceneManager.Models.Profile.startupScene","name":"startupScene","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_startupScene","commentId":"P:AdvancedSceneManager.Models.Profile.startupScene","fullName":"AdvancedSceneManager.Models.Profile.startupScene","nameWithType":"Profile.startupScene"},{"uid":"AdvancedSceneManager.Models.Profile.startupLoadingScreen","name":"startupLoadingScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_startupLoadingScreen","commentId":"P:AdvancedSceneManager.Models.Profile.startupLoadingScreen","fullName":"AdvancedSceneManager.Models.Profile.startupLoadingScreen","nameWithType":"Profile.startupLoadingScreen"},{"uid":"AdvancedSceneManager.Models.Profile.loadingScreen","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_loadingScreen","commentId":"P:AdvancedSceneManager.Models.Profile.loadingScreen","fullName":"AdvancedSceneManager.Models.Profile.loadingScreen","nameWithType":"Profile.loadingScreen"},{"uid":"AdvancedSceneManager.Models.Profile.splashScreen","name":"splashScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_splashScreen","commentId":"P:AdvancedSceneManager.Models.Profile.splashScreen","fullName":"AdvancedSceneManager.Models.Profile.splashScreen","nameWithType":"Profile.splashScreen"},{"uid":"AdvancedSceneManager.Models.Profile.useDefaultPauseScreen","name":"useDefaultPauseScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_useDefaultPauseScreen","commentId":"P:AdvancedSceneManager.Models.Profile.useDefaultPauseScreen","fullName":"AdvancedSceneManager.Models.Profile.useDefaultPauseScreen","nameWithType":"Profile.useDefaultPauseScreen"},{"uid":"AdvancedSceneManager.Models.Profile.includeFadeLoadingScene","name":"includeFadeLoadingScene","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_includeFadeLoadingScene","commentId":"P:AdvancedSceneManager.Models.Profile.includeFadeLoadingScene","fullName":"AdvancedSceneManager.Models.Profile.includeFadeLoadingScene","nameWithType":"Profile.includeFadeLoadingScene"},{"uid":"AdvancedSceneManager.Models.Profile.backgroundLoadingPriority","name":"backgroundLoadingPriority","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_backgroundLoadingPriority","commentId":"P:AdvancedSceneManager.Models.Profile.backgroundLoadingPriority","fullName":"AdvancedSceneManager.Models.Profile.backgroundLoadingPriority","nameWithType":"Profile.backgroundLoadingPriority"},{"uid":"AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority","name":"enableChangingBackgroundLoadingPriority","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_enableChangingBackgroundLoadingPriority","commentId":"P:AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority","fullName":"AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority","nameWithType":"Profile.enableChangingBackgroundLoadingPriority"},{"uid":"AdvancedSceneManager.Models.Profile.createCameraDuringStartup","name":"createCameraDuringStartup","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_createCameraDuringStartup","commentId":"P:AdvancedSceneManager.Models.Profile.createCameraDuringStartup","fullName":"AdvancedSceneManager.Models.Profile.createCameraDuringStartup","nameWithType":"Profile.createCameraDuringStartup"},{"uid":"AdvancedSceneManager.Models.Profile.tagDefinitions","name":"tagDefinitions","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_tagDefinitions","commentId":"F:AdvancedSceneManager.Models.Profile.tagDefinitions","fullName":"AdvancedSceneManager.Models.Profile.tagDefinitions","nameWithType":"Profile.tagDefinitions"},{"uid":"AdvancedSceneManager.Models.Profile.dynamicCollectionPaths","name":"dynamicCollectionPaths","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_dynamicCollectionPaths","commentId":"P:AdvancedSceneManager.Models.Profile.dynamicCollectionPaths","fullName":"AdvancedSceneManager.Models.Profile.dynamicCollectionPaths","nameWithType":"Profile.dynamicCollectionPaths"},{"uid":"AdvancedSceneManager.Models.Profile.blacklist","name":"blacklist","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_blacklist","commentId":"P:AdvancedSceneManager.Models.Profile.blacklist","fullName":"AdvancedSceneManager.Models.Profile.blacklist","nameWithType":"Profile.blacklist"},{"uid":"AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection)","name":"Order(SceneCollection)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Order_AdvancedSceneManager_Models_SceneCollection_","commentId":"M:AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection)","fullName":"AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection)","nameWithType":"Profile.Order(SceneCollection)"},{"uid":"AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32})","name":"Order(SceneCollection, Nullable<Int32>)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Order_AdvancedSceneManager_Models_SceneCollection_System_Nullable_System_Int32__","commentId":"M:AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection,System.Nullable{System.Int32})","name.vb":"Order(SceneCollection, Nullable(Of Int32))","fullName":"AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection, System.Nullable<System.Int32>)","fullName.vb":"AdvancedSceneManager.Models.Profile.Order(AdvancedSceneManager.Models.SceneCollection, System.Nullable(Of System.Int32))","nameWithType":"Profile.Order(SceneCollection, Nullable<Int32>)","nameWithType.vb":"Profile.Order(SceneCollection, Nullable(Of Int32))"},{"uid":"AdvancedSceneManager.Models.Profile.dynamicCollections","name":"dynamicCollections","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_dynamicCollections","commentId":"P:AdvancedSceneManager.Models.Profile.dynamicCollections","fullName":"AdvancedSceneManager.Models.Profile.dynamicCollections","nameWithType":"Profile.dynamicCollections"},{"uid":"AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.Scene,System.String,System.Boolean)","name":"Add(Scene, String, Boolean)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Add_AdvancedSceneManager_Models_Scene_System_String_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.Scene,System.String,System.Boolean)","fullName":"AdvancedSceneManager.Models.Profile.Add(AdvancedSceneManager.Models.Scene, System.String, System.Boolean)","nameWithType":"Profile.Add(Scene, String, Boolean)"},{"uid":"AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.Scene,System.String,System.Boolean)","name":"Remove(Scene, String, Boolean)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Remove_AdvancedSceneManager_Models_Scene_System_String_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.Scene,System.String,System.Boolean)","fullName":"AdvancedSceneManager.Models.Profile.Remove(AdvancedSceneManager.Models.Scene, System.String, System.Boolean)","nameWithType":"Profile.Remove(Scene, String, Boolean)"},{"uid":"AdvancedSceneManager.Models.Profile.Clear(System.String,System.Boolean,System.Boolean)","name":"Clear(String, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Clear_System_String_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Profile.Clear(System.String,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Models.Profile.Clear(System.String, System.Boolean, System.Boolean)","nameWithType":"Profile.Clear(String, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Models.Profile.IsSet(System.String,System.String)","name":"IsSet(String, String)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_IsSet_System_String_System_String_","commentId":"M:AdvancedSceneManager.Models.Profile.IsSet(System.String,System.String)","fullName":"AdvancedSceneManager.Models.Profile.IsSet(System.String, System.String)","nameWithType":"Profile.IsSet(String, String)"},{"uid":"AdvancedSceneManager.Models.Profile.IsSet(System.String,System.Boolean)","name":"IsSet(String, Boolean)","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_IsSet_System_String_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Profile.IsSet(System.String,System.Boolean)","fullName":"AdvancedSceneManager.Models.Profile.IsSet(System.String, System.Boolean)","nameWithType":"Profile.IsSet(String, Boolean)"},{"uid":"AdvancedSceneManager.Models.Profile.Delete","name":"Delete()","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Delete","commentId":"M:AdvancedSceneManager.Models.Profile.Delete","fullName":"AdvancedSceneManager.Models.Profile.Delete()","nameWithType":"Profile.Delete()"},{"uid":"AdvancedSceneManager.Models.Profile.FindAll*","name":"FindAll","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_FindAll_","commentId":"Overload:AdvancedSceneManager.Models.Profile.FindAll","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.FindAll","nameWithType":"Profile.FindAll"},{"uid":"AdvancedSceneManager.Models.Profile.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Find_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Find","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Find","nameWithType":"Profile.Find"},{"uid":"AdvancedSceneManager.Models.Profile.name*","name":"name","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_name_","commentId":"Overload:AdvancedSceneManager.Models.Profile.name","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.name","nameWithType":"Profile.name"},{"uid":"AdvancedSceneManager.Models.Profile.MarkAsDirty*","name":"MarkAsDirty","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_MarkAsDirty_","commentId":"Overload:AdvancedSceneManager.Models.Profile.MarkAsDirty","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.MarkAsDirty","nameWithType":"Profile.MarkAsDirty"},{"uid":"AdvancedSceneManager.Models.Profile.current*","name":"current","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_current_","commentId":"Overload:AdvancedSceneManager.Models.Profile.current","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.current","nameWithType":"Profile.current"},{"uid":"AdvancedSceneManager.Models.Profile.collections*","name":"collections","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_collections_","commentId":"Overload:AdvancedSceneManager.Models.Profile.collections","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.collections","nameWithType":"Profile.collections"},{"uid":"AdvancedSceneManager.Models.Profile.scenes*","name":"scenes","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_scenes_","commentId":"Overload:AdvancedSceneManager.Models.Profile.scenes","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.scenes","nameWithType":"Profile.scenes"},{"uid":"AdvancedSceneManager.Models.Profile.scenePaths*","name":"scenePaths","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_scenePaths_","commentId":"Overload:AdvancedSceneManager.Models.Profile.scenePaths","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.scenePaths","nameWithType":"Profile.scenePaths"},{"uid":"AdvancedSceneManager.Models.Profile.StartupCollections*","name":"StartupCollections","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_StartupCollections_","commentId":"Overload:AdvancedSceneManager.Models.Profile.StartupCollections","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.StartupCollections","nameWithType":"Profile.StartupCollections"},{"uid":"AdvancedSceneManager.Models.Profile.CreateCollection*","name":"CreateCollection","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_CreateCollection_","commentId":"Overload:AdvancedSceneManager.Models.Profile.CreateCollection","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.CreateCollection","nameWithType":"Profile.CreateCollection"},{"uid":"AdvancedSceneManager.Models.Profile.Add*","name":"Add","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Add_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Add","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Add","nameWithType":"Profile.Add"},{"uid":"AdvancedSceneManager.Models.Profile.Remove*","name":"Remove","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Remove_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Remove","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Remove","nameWithType":"Profile.Remove"},{"uid":"AdvancedSceneManager.Models.Profile.startupScene*","name":"startupScene","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_startupScene_","commentId":"Overload:AdvancedSceneManager.Models.Profile.startupScene","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.startupScene","nameWithType":"Profile.startupScene"},{"uid":"AdvancedSceneManager.Models.Profile.startupLoadingScreen*","name":"startupLoadingScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_startupLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Models.Profile.startupLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.startupLoadingScreen","nameWithType":"Profile.startupLoadingScreen"},{"uid":"AdvancedSceneManager.Models.Profile.loadingScreen*","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_loadingScreen_","commentId":"Overload:AdvancedSceneManager.Models.Profile.loadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.loadingScreen","nameWithType":"Profile.loadingScreen"},{"uid":"AdvancedSceneManager.Models.Profile.splashScreen*","name":"splashScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_splashScreen_","commentId":"Overload:AdvancedSceneManager.Models.Profile.splashScreen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.splashScreen","nameWithType":"Profile.splashScreen"},{"uid":"AdvancedSceneManager.Models.Profile.useDefaultPauseScreen*","name":"useDefaultPauseScreen","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_useDefaultPauseScreen_","commentId":"Overload:AdvancedSceneManager.Models.Profile.useDefaultPauseScreen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.useDefaultPauseScreen","nameWithType":"Profile.useDefaultPauseScreen"},{"uid":"AdvancedSceneManager.Models.Profile.includeFadeLoadingScene*","name":"includeFadeLoadingScene","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_includeFadeLoadingScene_","commentId":"Overload:AdvancedSceneManager.Models.Profile.includeFadeLoadingScene","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.includeFadeLoadingScene","nameWithType":"Profile.includeFadeLoadingScene"},{"uid":"AdvancedSceneManager.Models.Profile.backgroundLoadingPriority*","name":"backgroundLoadingPriority","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_backgroundLoadingPriority_","commentId":"Overload:AdvancedSceneManager.Models.Profile.backgroundLoadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.backgroundLoadingPriority","nameWithType":"Profile.backgroundLoadingPriority"},{"uid":"AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority*","name":"enableChangingBackgroundLoadingPriority","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_enableChangingBackgroundLoadingPriority_","commentId":"Overload:AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.enableChangingBackgroundLoadingPriority","nameWithType":"Profile.enableChangingBackgroundLoadingPriority"},{"uid":"AdvancedSceneManager.Models.Profile.createCameraDuringStartup*","name":"createCameraDuringStartup","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_createCameraDuringStartup_","commentId":"Overload:AdvancedSceneManager.Models.Profile.createCameraDuringStartup","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.createCameraDuringStartup","nameWithType":"Profile.createCameraDuringStartup"},{"uid":"AdvancedSceneManager.Models.Profile.dynamicCollectionPaths*","name":"dynamicCollectionPaths","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_dynamicCollectionPaths_","commentId":"Overload:AdvancedSceneManager.Models.Profile.dynamicCollectionPaths","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.dynamicCollectionPaths","nameWithType":"Profile.dynamicCollectionPaths"},{"uid":"AdvancedSceneManager.Models.Profile.blacklist*","name":"blacklist","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_blacklist_","commentId":"Overload:AdvancedSceneManager.Models.Profile.blacklist","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.blacklist","nameWithType":"Profile.blacklist"},{"uid":"AdvancedSceneManager.Models.Profile.Order*","name":"Order","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Order_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Order","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Order","nameWithType":"Profile.Order"},{"uid":"AdvancedSceneManager.Models.Profile.dynamicCollections*","name":"dynamicCollections","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_dynamicCollections_","commentId":"Overload:AdvancedSceneManager.Models.Profile.dynamicCollections","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.dynamicCollections","nameWithType":"Profile.dynamicCollections"},{"uid":"AdvancedSceneManager.Models.Profile.Clear*","name":"Clear","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Clear_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Clear","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Clear","nameWithType":"Profile.Clear"},{"uid":"AdvancedSceneManager.Models.Profile.IsSet*","name":"IsSet","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_IsSet_","commentId":"Overload:AdvancedSceneManager.Models.Profile.IsSet","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.IsSet","nameWithType":"Profile.IsSet"},{"uid":"AdvancedSceneManager.Models.Profile.Delete*","name":"Delete","href":"~/api/AdvancedSceneManager.Models.Profile.yml#AdvancedSceneManager_Models_Profile_Delete_","commentId":"Overload:AdvancedSceneManager.Models.Profile.Delete","isSpec":"True","fullName":"AdvancedSceneManager.Models.Profile.Delete","nameWithType":"Profile.Delete"}],"api/AdvancedSceneManager.Models.Scene.yml":[{"uid":"AdvancedSceneManager.Models.Scene","name":"Scene","href":"~/api/AdvancedSceneManager.Models.Scene.yml","commentId":"T:AdvancedSceneManager.Models.Scene","fullName":"AdvancedSceneManager.Models.Scene","nameWithType":"Scene"},{"uid":"AdvancedSceneManager.Models.Scene.PropertyChanged","name":"PropertyChanged","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_PropertyChanged","commentId":"E:AdvancedSceneManager.Models.Scene.PropertyChanged","fullName":"AdvancedSceneManager.Models.Scene.PropertyChanged","nameWithType":"Scene.PropertyChanged"},{"uid":"AdvancedSceneManager.Models.Scene.OnPropertyChanged","name":"OnPropertyChanged()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OnPropertyChanged","commentId":"M:AdvancedSceneManager.Models.Scene.OnPropertyChanged","fullName":"AdvancedSceneManager.Models.Scene.OnPropertyChanged()","nameWithType":"Scene.OnPropertyChanged()"},{"uid":"AdvancedSceneManager.Models.Scene.name","name":"name","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_name","commentId":"P:AdvancedSceneManager.Models.Scene.name","fullName":"AdvancedSceneManager.Models.Scene.name","nameWithType":"Scene.name"},{"uid":"AdvancedSceneManager.Models.Scene.path","name":"path","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_path","commentId":"P:AdvancedSceneManager.Models.Scene.path","fullName":"AdvancedSceneManager.Models.Scene.path","nameWithType":"Scene.path"},{"uid":"AdvancedSceneManager.Models.Scene.assetID","name":"assetID","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_assetID","commentId":"P:AdvancedSceneManager.Models.Scene.assetID","fullName":"AdvancedSceneManager.Models.Scene.assetID","nameWithType":"Scene.assetID"},{"uid":"AdvancedSceneManager.Models.Scene.isIncluded","name":"isIncluded","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_isIncluded","commentId":"P:AdvancedSceneManager.Models.Scene.isIncluded","fullName":"AdvancedSceneManager.Models.Scene.isIncluded","nameWithType":"Scene.isIncluded"},{"uid":"AdvancedSceneManager.Models.Scene.isActive","name":"isActive","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_isActive","commentId":"P:AdvancedSceneManager.Models.Scene.isActive","fullName":"AdvancedSceneManager.Models.Scene.isActive","nameWithType":"Scene.isActive"},{"uid":"AdvancedSceneManager.Models.Scene.SetActiveScene","name":"SetActiveScene()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_SetActiveScene","commentId":"M:AdvancedSceneManager.Models.Scene.SetActiveScene","fullName":"AdvancedSceneManager.Models.Scene.SetActiveScene()","nameWithType":"Scene.SetActiveScene()"},{"uid":"AdvancedSceneManager.Models.Scene.IsOpen","name":"IsOpen()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_IsOpen","commentId":"M:AdvancedSceneManager.Models.Scene.IsOpen","fullName":"AdvancedSceneManager.Models.Scene.IsOpen()","nameWithType":"Scene.IsOpen()"},{"uid":"AdvancedSceneManager.Models.Scene.Open","name":"Open()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Open","commentId":"M:AdvancedSceneManager.Models.Scene.Open","fullName":"AdvancedSceneManager.Models.Scene.Open()","nameWithType":"Scene.Open()"},{"uid":"AdvancedSceneManager.Models.Scene.OpenSingle","name":"OpenSingle()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenSingle","commentId":"M:AdvancedSceneManager.Models.Scene.OpenSingle","fullName":"AdvancedSceneManager.Models.Scene.OpenSingle()","nameWithType":"Scene.OpenSingle()"},{"uid":"AdvancedSceneManager.Models.Scene.Reopen","name":"Reopen()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Reopen","commentId":"M:AdvancedSceneManager.Models.Scene.Reopen","fullName":"AdvancedSceneManager.Models.Scene.Reopen()","nameWithType":"Scene.Reopen()"},{"uid":"AdvancedSceneManager.Models.Scene.Toggle","name":"Toggle()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Toggle","commentId":"M:AdvancedSceneManager.Models.Scene.Toggle","fullName":"AdvancedSceneManager.Models.Scene.Toggle()","nameWithType":"Scene.Toggle()"},{"uid":"AdvancedSceneManager.Models.Scene.Toggle(System.Boolean)","name":"Toggle(Boolean)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Toggle_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Scene.Toggle(System.Boolean)","fullName":"AdvancedSceneManager.Models.Scene.Toggle(System.Boolean)","nameWithType":"Scene.Toggle(Boolean)"},{"uid":"AdvancedSceneManager.Models.Scene.Close","name":"Close()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Close","commentId":"M:AdvancedSceneManager.Models.Scene.Close","fullName":"AdvancedSceneManager.Models.Scene.Close()","nameWithType":"Scene.Close()"},{"uid":"AdvancedSceneManager.Models.Scene.Preload","name":"Preload()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Preload","commentId":"M:AdvancedSceneManager.Models.Scene.Preload","fullName":"AdvancedSceneManager.Models.Scene.Preload()","nameWithType":"Scene.Preload()"},{"uid":"AdvancedSceneManager.Models.Scene.OpenEvent","name":"OpenEvent()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenEvent","commentId":"M:AdvancedSceneManager.Models.Scene.OpenEvent","fullName":"AdvancedSceneManager.Models.Scene.OpenEvent()","nameWithType":"Scene.OpenEvent()"},{"uid":"AdvancedSceneManager.Models.Scene.OpenSingleEvent","name":"OpenSingleEvent()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenSingleEvent","commentId":"M:AdvancedSceneManager.Models.Scene.OpenSingleEvent","fullName":"AdvancedSceneManager.Models.Scene.OpenSingleEvent()","nameWithType":"Scene.OpenSingleEvent()"},{"uid":"AdvancedSceneManager.Models.Scene.ReopenEvent","name":"ReopenEvent()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_ReopenEvent","commentId":"M:AdvancedSceneManager.Models.Scene.ReopenEvent","fullName":"AdvancedSceneManager.Models.Scene.ReopenEvent()","nameWithType":"Scene.ReopenEvent()"},{"uid":"AdvancedSceneManager.Models.Scene.ToggleEvent","name":"ToggleEvent()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_ToggleEvent","commentId":"M:AdvancedSceneManager.Models.Scene.ToggleEvent","fullName":"AdvancedSceneManager.Models.Scene.ToggleEvent()","nameWithType":"Scene.ToggleEvent()"},{"uid":"AdvancedSceneManager.Models.Scene.ToggleEvent(System.Boolean)","name":"ToggleEvent(Boolean)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_ToggleEvent_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Scene.ToggleEvent(System.Boolean)","fullName":"AdvancedSceneManager.Models.Scene.ToggleEvent(System.Boolean)","nameWithType":"Scene.ToggleEvent(Boolean)"},{"uid":"AdvancedSceneManager.Models.Scene.CloseEvent","name":"CloseEvent()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_CloseEvent","commentId":"M:AdvancedSceneManager.Models.Scene.CloseEvent","fullName":"AdvancedSceneManager.Models.Scene.CloseEvent()","nameWithType":"Scene.CloseEvent()"},{"uid":"AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent(AdvancedSceneManager.Models.Scene)","name":"OpenWithLoadingScreenEvent(Scene)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenWithLoadingScreenEvent_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent(AdvancedSceneManager.Models.Scene)","nameWithType":"Scene.OpenWithLoadingScreenEvent(Scene)"},{"uid":"AdvancedSceneManager.Models.Scene.GetOpenSceneInfo","name":"GetOpenSceneInfo()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetOpenSceneInfo","commentId":"M:AdvancedSceneManager.Models.Scene.GetOpenSceneInfo","fullName":"AdvancedSceneManager.Models.Scene.GetOpenSceneInfo()","nameWithType":"Scene.GetOpenSceneInfo()"},{"uid":"AdvancedSceneManager.Models.Scene.FindCollections(System.Boolean)","name":"FindCollections(Boolean)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindCollections_System_Boolean_","commentId":"M:AdvancedSceneManager.Models.Scene.FindCollections(System.Boolean)","fullName":"AdvancedSceneManager.Models.Scene.FindCollections(System.Boolean)","nameWithType":"Scene.FindCollections(Boolean)"},{"uid":"AdvancedSceneManager.Models.Scene.FindCollections(AdvancedSceneManager.Models.Profile)","name":"FindCollections(Profile)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindCollections_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Models.Scene.FindCollections(AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Models.Scene.FindCollections(AdvancedSceneManager.Models.Profile)","nameWithType":"Scene.FindCollections(Profile)"},{"uid":"AdvancedSceneManager.Models.Scene.GetRootGameObjects","name":"GetRootGameObjects()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetRootGameObjects","commentId":"M:AdvancedSceneManager.Models.Scene.GetRootGameObjects","fullName":"AdvancedSceneManager.Models.Scene.GetRootGameObjects()","nameWithType":"Scene.GetRootGameObjects()"},{"uid":"AdvancedSceneManager.Models.Scene.FindObject``1","name":"FindObject<T>()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindObject__1","commentId":"M:AdvancedSceneManager.Models.Scene.FindObject``1","name.vb":"FindObject(Of T)()","fullName":"AdvancedSceneManager.Models.Scene.FindObject<T>()","fullName.vb":"AdvancedSceneManager.Models.Scene.FindObject(Of T)()","nameWithType":"Scene.FindObject<T>()","nameWithType.vb":"Scene.FindObject(Of T)()"},{"uid":"AdvancedSceneManager.Models.Scene.FindObjects``1","name":"FindObjects<T>()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindObjects__1","commentId":"M:AdvancedSceneManager.Models.Scene.FindObjects``1","name.vb":"FindObjects(Of T)()","fullName":"AdvancedSceneManager.Models.Scene.FindObjects<T>()","fullName.vb":"AdvancedSceneManager.Models.Scene.FindObjects(Of T)()","nameWithType":"Scene.FindObjects<T>()","nameWithType.vb":"Scene.FindObjects(Of T)()"},{"uid":"AdvancedSceneManager.Models.Scene.Find(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name":"Find(String, SceneCollection, Profile)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Find_System_String_AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Models.Scene.Find(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Models.Scene.Find(System.String, AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","nameWithType":"Scene.Find(String, SceneCollection, Profile)"},{"uid":"AdvancedSceneManager.Models.Scene.FindAll(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","name":"FindAll(String, SceneCollection, Profile)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindAll_System_String_AdvancedSceneManager_Models_SceneCollection_AdvancedSceneManager_Models_Profile_","commentId":"M:AdvancedSceneManager.Models.Scene.FindAll(System.String,AdvancedSceneManager.Models.SceneCollection,AdvancedSceneManager.Models.Profile)","fullName":"AdvancedSceneManager.Models.Scene.FindAll(System.String, AdvancedSceneManager.Models.SceneCollection, AdvancedSceneManager.Models.Profile)","nameWithType":"Scene.FindAll(String, SceneCollection, Profile)"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(System.Object)","name":"Equals(Object)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_System_Object_","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(System.Object)","fullName":"AdvancedSceneManager.Models.Scene.Equals(System.Object)","nameWithType":"Scene.Equals(Object)"},{"uid":"AdvancedSceneManager.Models.Scene.GetHashCode","name":"GetHashCode()","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetHashCode","commentId":"M:AdvancedSceneManager.Models.Scene.GetHashCode","fullName":"AdvancedSceneManager.Models.Scene.GetHashCode()","nameWithType":"Scene.GetHashCode()"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Models.Scene)","name":"Equals(Scene)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Models.Scene)","nameWithType":"Scene.Equals(Scene)"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","name":"Equals(OpenSceneInfo)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_AdvancedSceneManager_Core_OpenSceneInfo_","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","fullName":"AdvancedSceneManager.Models.Scene.Equals(AdvancedSceneManager.Core.OpenSceneInfo)","nameWithType":"Scene.Equals(OpenSceneInfo)"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(UnityEngine.SceneManagement.Scene)","name":"Equals(Scene)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Models.Scene.Equals(UnityEngine.SceneManagement.Scene)","nameWithType":"Scene.Equals(Scene)"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(System.Nullable{UnityEngine.SceneManagement.Scene})","name":"Equals(Nullable<Scene>)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_System_Nullable_UnityEngine_SceneManagement_Scene__","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(System.Nullable{UnityEngine.SceneManagement.Scene})","name.vb":"Equals(Nullable(Of Scene))","fullName":"AdvancedSceneManager.Models.Scene.Equals(System.Nullable<UnityEngine.SceneManagement.Scene>)","fullName.vb":"AdvancedSceneManager.Models.Scene.Equals(System.Nullable(Of UnityEngine.SceneManagement.Scene))","nameWithType":"Scene.Equals(Nullable<Scene>)","nameWithType.vb":"Scene.Equals(Nullable(Of Scene))"},{"uid":"AdvancedSceneManager.Models.Scene.Equals(UnityEditor.SceneAsset)","name":"Equals(SceneAsset)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_UnityEditor_SceneAsset_","commentId":"M:AdvancedSceneManager.Models.Scene.Equals(UnityEditor.SceneAsset)","fullName":"AdvancedSceneManager.Models.Scene.Equals(UnityEditor.SceneAsset)","nameWithType":"Scene.Equals(SceneAsset)"},{"uid":"AdvancedSceneManager.Models.Scene.OnOpen(System.Int32,System.Int32)","name":"OnOpen(Int32, Int32)","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OnOpen_System_Int32_System_Int32_","commentId":"M:AdvancedSceneManager.Models.Scene.OnOpen(System.Int32,System.Int32)","fullName":"AdvancedSceneManager.Models.Scene.OnOpen(System.Int32, System.Int32)","nameWithType":"Scene.OnOpen(Int32, Int32)"},{"uid":"AdvancedSceneManager.Models.Scene.OnPropertyChanged*","name":"OnPropertyChanged","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OnPropertyChanged_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OnPropertyChanged","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OnPropertyChanged","nameWithType":"Scene.OnPropertyChanged"},{"uid":"AdvancedSceneManager.Models.Scene.name*","name":"name","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_name_","commentId":"Overload:AdvancedSceneManager.Models.Scene.name","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.name","nameWithType":"Scene.name"},{"uid":"AdvancedSceneManager.Models.Scene.path*","name":"path","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_path_","commentId":"Overload:AdvancedSceneManager.Models.Scene.path","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.path","nameWithType":"Scene.path"},{"uid":"AdvancedSceneManager.Models.Scene.assetID*","name":"assetID","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_assetID_","commentId":"Overload:AdvancedSceneManager.Models.Scene.assetID","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.assetID","nameWithType":"Scene.assetID"},{"uid":"AdvancedSceneManager.Models.Scene.isIncluded*","name":"isIncluded","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_isIncluded_","commentId":"Overload:AdvancedSceneManager.Models.Scene.isIncluded","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.isIncluded","nameWithType":"Scene.isIncluded"},{"uid":"AdvancedSceneManager.Models.Scene.isActive*","name":"isActive","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_isActive_","commentId":"Overload:AdvancedSceneManager.Models.Scene.isActive","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.isActive","nameWithType":"Scene.isActive"},{"uid":"AdvancedSceneManager.Models.Scene.SetActiveScene*","name":"SetActiveScene","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_SetActiveScene_","commentId":"Overload:AdvancedSceneManager.Models.Scene.SetActiveScene","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.SetActiveScene","nameWithType":"Scene.SetActiveScene"},{"uid":"AdvancedSceneManager.Models.Scene.IsOpen*","name":"IsOpen","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_IsOpen_","commentId":"Overload:AdvancedSceneManager.Models.Scene.IsOpen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.IsOpen","nameWithType":"Scene.IsOpen"},{"uid":"AdvancedSceneManager.Models.Scene.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Open_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Open","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Open","nameWithType":"Scene.Open"},{"uid":"AdvancedSceneManager.Models.Scene.OpenSingle*","name":"OpenSingle","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenSingle_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OpenSingle","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OpenSingle","nameWithType":"Scene.OpenSingle"},{"uid":"AdvancedSceneManager.Models.Scene.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Reopen_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Reopen","nameWithType":"Scene.Reopen"},{"uid":"AdvancedSceneManager.Models.Scene.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Toggle_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Toggle","nameWithType":"Scene.Toggle"},{"uid":"AdvancedSceneManager.Models.Scene.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Close_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Close","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Close","nameWithType":"Scene.Close"},{"uid":"AdvancedSceneManager.Models.Scene.Preload*","name":"Preload","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Preload_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Preload","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Preload","nameWithType":"Scene.Preload"},{"uid":"AdvancedSceneManager.Models.Scene.OpenEvent*","name":"OpenEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OpenEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OpenEvent","nameWithType":"Scene.OpenEvent"},{"uid":"AdvancedSceneManager.Models.Scene.OpenSingleEvent*","name":"OpenSingleEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenSingleEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OpenSingleEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OpenSingleEvent","nameWithType":"Scene.OpenSingleEvent"},{"uid":"AdvancedSceneManager.Models.Scene.ReopenEvent*","name":"ReopenEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_ReopenEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.ReopenEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.ReopenEvent","nameWithType":"Scene.ReopenEvent"},{"uid":"AdvancedSceneManager.Models.Scene.ToggleEvent*","name":"ToggleEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_ToggleEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.ToggleEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.ToggleEvent","nameWithType":"Scene.ToggleEvent"},{"uid":"AdvancedSceneManager.Models.Scene.CloseEvent*","name":"CloseEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_CloseEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.CloseEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.CloseEvent","nameWithType":"Scene.CloseEvent"},{"uid":"AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent*","name":"OpenWithLoadingScreenEvent","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OpenWithLoadingScreenEvent_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OpenWithLoadingScreenEvent","nameWithType":"Scene.OpenWithLoadingScreenEvent"},{"uid":"AdvancedSceneManager.Models.Scene.GetOpenSceneInfo*","name":"GetOpenSceneInfo","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetOpenSceneInfo_","commentId":"Overload:AdvancedSceneManager.Models.Scene.GetOpenSceneInfo","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.GetOpenSceneInfo","nameWithType":"Scene.GetOpenSceneInfo"},{"uid":"AdvancedSceneManager.Models.Scene.FindCollections*","name":"FindCollections","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindCollections_","commentId":"Overload:AdvancedSceneManager.Models.Scene.FindCollections","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.FindCollections","nameWithType":"Scene.FindCollections"},{"uid":"AdvancedSceneManager.Models.Scene.GetRootGameObjects*","name":"GetRootGameObjects","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetRootGameObjects_","commentId":"Overload:AdvancedSceneManager.Models.Scene.GetRootGameObjects","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.GetRootGameObjects","nameWithType":"Scene.GetRootGameObjects"},{"uid":"AdvancedSceneManager.Models.Scene.FindObject*","name":"FindObject","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindObject_","commentId":"Overload:AdvancedSceneManager.Models.Scene.FindObject","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.FindObject","nameWithType":"Scene.FindObject"},{"uid":"AdvancedSceneManager.Models.Scene.FindObjects*","name":"FindObjects","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindObjects_","commentId":"Overload:AdvancedSceneManager.Models.Scene.FindObjects","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.FindObjects","nameWithType":"Scene.FindObjects"},{"uid":"AdvancedSceneManager.Models.Scene.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Find_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Find","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Find","nameWithType":"Scene.Find"},{"uid":"AdvancedSceneManager.Models.Scene.FindAll*","name":"FindAll","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_FindAll_","commentId":"Overload:AdvancedSceneManager.Models.Scene.FindAll","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.FindAll","nameWithType":"Scene.FindAll"},{"uid":"AdvancedSceneManager.Models.Scene.Equals*","name":"Equals","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_Equals_","commentId":"Overload:AdvancedSceneManager.Models.Scene.Equals","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.Equals","nameWithType":"Scene.Equals"},{"uid":"AdvancedSceneManager.Models.Scene.GetHashCode*","name":"GetHashCode","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_GetHashCode_","commentId":"Overload:AdvancedSceneManager.Models.Scene.GetHashCode","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.GetHashCode","nameWithType":"Scene.GetHashCode"},{"uid":"AdvancedSceneManager.Models.Scene.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Models.Scene.yml#AdvancedSceneManager_Models_Scene_OnOpen_","commentId":"Overload:AdvancedSceneManager.Models.Scene.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Models.Scene.OnOpen","nameWithType":"Scene.OnOpen"}],"api/AdvancedSceneManager.Utility.PauseScreenUtility.yml":[{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility","name":"PauseScreenUtility","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml","commentId":"T:AdvancedSceneManager.Utility.PauseScreenUtility","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility","nameWithType":"PauseScreenUtility"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.isOpen","name":"isOpen","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_isOpen","commentId":"P:AdvancedSceneManager.Utility.PauseScreenUtility.isOpen","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.isOpen","nameWithType":"PauseScreenUtility.isOpen"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey","name":"ListenForKey()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_ListenForKey","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey()","nameWithType":"PauseScreenUtility.ListenForKey()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.StopListening","name":"StopListening()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_StopListening","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.StopListening","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.StopListening()","nameWithType":"PauseScreenUtility.StopListening()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Show","name":"Show()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Show","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Show","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Show()","nameWithType":"PauseScreenUtility.Show()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Hide(System.Boolean)","name":"Hide(Boolean)","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Hide_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Hide(System.Boolean)","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Hide(System.Boolean)","nameWithType":"PauseScreenUtility.Hide(Boolean)"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Toggle","name":"Toggle()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Toggle","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Toggle","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Toggle()","nameWithType":"PauseScreenUtility.Toggle()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.resume","name":"resume","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_resume","commentId":"F:AdvancedSceneManager.Utility.PauseScreenUtility.resume","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.resume","nameWithType":"PauseScreenUtility.resume"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.restartCollection","name":"restartCollection","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_restartCollection","commentId":"F:AdvancedSceneManager.Utility.PauseScreenUtility.restartCollection","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.restartCollection","nameWithType":"PauseScreenUtility.restartCollection"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.restartGame","name":"restartGame","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_restartGame","commentId":"F:AdvancedSceneManager.Utility.PauseScreenUtility.restartGame","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.restartGame","nameWithType":"PauseScreenUtility.restartGame"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.quit","name":"quit","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_quit","commentId":"F:AdvancedSceneManager.Utility.PauseScreenUtility.quit","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.quit","nameWithType":"PauseScreenUtility.quit"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.canvasGroup","name":"canvasGroup","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_canvasGroup","commentId":"F:AdvancedSceneManager.Utility.PauseScreenUtility.canvasGroup","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.canvasGroup","nameWithType":"PauseScreenUtility.canvasGroup"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Begin","name":"Begin()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Begin","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Begin","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Begin()","nameWithType":"PauseScreenUtility.Begin()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.End","name":"End()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_End","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.End","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.End()","nameWithType":"PauseScreenUtility.End()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection","name":"RestartCollection()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_RestartCollection","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection()","nameWithType":"PauseScreenUtility.RestartCollection()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame","name":"RestartGame()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_RestartGame","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame()","nameWithType":"PauseScreenUtility.RestartGame()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Resume","name":"Resume()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Resume","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Resume","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Resume()","nameWithType":"PauseScreenUtility.Resume()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Quit","name":"Quit()","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Quit","commentId":"M:AdvancedSceneManager.Utility.PauseScreenUtility.Quit","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Quit()","nameWithType":"PauseScreenUtility.Quit()"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.isOpen*","name":"isOpen","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_isOpen_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.isOpen","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.isOpen","nameWithType":"PauseScreenUtility.isOpen"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey*","name":"ListenForKey","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_ListenForKey_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.ListenForKey","nameWithType":"PauseScreenUtility.ListenForKey"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.StopListening*","name":"StopListening","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_StopListening_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.StopListening","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.StopListening","nameWithType":"PauseScreenUtility.StopListening"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Show*","name":"Show","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Show_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Show","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Show","nameWithType":"PauseScreenUtility.Show"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Hide*","name":"Hide","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Hide_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Hide","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Hide","nameWithType":"PauseScreenUtility.Hide"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Toggle*","name":"Toggle","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Toggle_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Toggle","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Toggle","nameWithType":"PauseScreenUtility.Toggle"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Begin*","name":"Begin","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Begin_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Begin","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Begin","nameWithType":"PauseScreenUtility.Begin"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.End*","name":"End","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_End_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.End","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.End","nameWithType":"PauseScreenUtility.End"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection*","name":"RestartCollection","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_RestartCollection_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartCollection","nameWithType":"PauseScreenUtility.RestartCollection"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame*","name":"RestartGame","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_RestartGame_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.RestartGame","nameWithType":"PauseScreenUtility.RestartGame"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Resume*","name":"Resume","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Resume_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Resume","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Resume","nameWithType":"PauseScreenUtility.Resume"},{"uid":"AdvancedSceneManager.Utility.PauseScreenUtility.Quit*","name":"Quit","href":"~/api/AdvancedSceneManager.Utility.PauseScreenUtility.yml#AdvancedSceneManager_Utility_PauseScreenUtility_Quit_","commentId":"Overload:AdvancedSceneManager.Utility.PauseScreenUtility.Quit","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PauseScreenUtility.Quit","nameWithType":"PauseScreenUtility.Quit"}],"api/AdvancedSceneManager.Utility.PersistentUtility.yml":[{"uid":"AdvancedSceneManager.Utility.PersistentUtility","name":"PersistentUtility","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml","commentId":"T:AdvancedSceneManager.Utility.PersistentUtility","fullName":"AdvancedSceneManager.Utility.PersistentUtility","nameWithType":"PersistentUtility"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.Set(UnityEngine.SceneManagement.Scene,AdvancedSceneManager.Models.SceneCloseBehavior)","name":"Set(Scene, SceneCloseBehavior)","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_Set_UnityEngine_SceneManagement_Scene_AdvancedSceneManager_Models_SceneCloseBehavior_","commentId":"M:AdvancedSceneManager.Utility.PersistentUtility.Set(UnityEngine.SceneManagement.Scene,AdvancedSceneManager.Models.SceneCloseBehavior)","fullName":"AdvancedSceneManager.Utility.PersistentUtility.Set(UnityEngine.SceneManagement.Scene, AdvancedSceneManager.Models.SceneCloseBehavior)","nameWithType":"PersistentUtility.Set(Scene, SceneCloseBehavior)"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.Unset(UnityEngine.SceneManagement.Scene)","name":"Unset(Scene)","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_Unset_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.PersistentUtility.Unset(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.PersistentUtility.Unset(UnityEngine.SceneManagement.Scene)","nameWithType":"PersistentUtility.Unset(Scene)"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.UnsetAll","name":"UnsetAll()","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_UnsetAll","commentId":"M:AdvancedSceneManager.Utility.PersistentUtility.UnsetAll","fullName":"AdvancedSceneManager.Utility.PersistentUtility.UnsetAll()","nameWithType":"PersistentUtility.UnsetAll()"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption(UnityEngine.SceneManagement.Scene)","name":"GetPersistentOption(Scene)","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_GetPersistentOption_UnityEngine_SceneManagement_Scene_","commentId":"M:AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption(UnityEngine.SceneManagement.Scene)","fullName":"AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption(UnityEngine.SceneManagement.Scene)","nameWithType":"PersistentUtility.GetPersistentOption(Scene)"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.Set*","name":"Set","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_Set_","commentId":"Overload:AdvancedSceneManager.Utility.PersistentUtility.Set","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PersistentUtility.Set","nameWithType":"PersistentUtility.Set"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.Unset*","name":"Unset","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_Unset_","commentId":"Overload:AdvancedSceneManager.Utility.PersistentUtility.Unset","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PersistentUtility.Unset","nameWithType":"PersistentUtility.Unset"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.UnsetAll*","name":"UnsetAll","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_UnsetAll_","commentId":"Overload:AdvancedSceneManager.Utility.PersistentUtility.UnsetAll","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PersistentUtility.UnsetAll","nameWithType":"PersistentUtility.UnsetAll"},{"uid":"AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption*","name":"GetPersistentOption","href":"~/api/AdvancedSceneManager.Utility.PersistentUtility.yml#AdvancedSceneManager_Utility_PersistentUtility_GetPersistentOption_","commentId":"Overload:AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PersistentUtility.GetPersistentOption","nameWithType":"PersistentUtility.GetPersistentOption"}],"api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml":[{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper","name":"PreloadedSceneHelper","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml","commentId":"T:AdvancedSceneManager.Utility.PreloadedSceneHelper","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper","nameWithType":"PreloadedSceneHelper"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,System.Boolean)","name":"PreloadedSceneHelper(OpenSceneInfo, Boolean)","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper__ctor_AdvancedSceneManager_Core_OpenSceneInfo_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.PreloadedSceneHelper.#ctor(AdvancedSceneManager.Core.OpenSceneInfo,System.Boolean)","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.PreloadedSceneHelper(AdvancedSceneManager.Core.OpenSceneInfo, System.Boolean)","nameWithType":"PreloadedSceneHelper.PreloadedSceneHelper(OpenSceneInfo, Boolean)"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.scene","name":"scene","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_scene","commentId":"P:AdvancedSceneManager.Utility.PreloadedSceneHelper.scene","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.scene","nameWithType":"PreloadedSceneHelper.scene"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded","name":"isStillPreloaded","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_isStillPreloaded","commentId":"P:AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded","nameWithType":"PreloadedSceneHelper.isStillPreloaded"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks","name":"hasRunCallbacks","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_hasRunCallbacks","commentId":"P:AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks","nameWithType":"PreloadedSceneHelper.hasRunCallbacks"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading","name":"FinishLoading()","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_FinishLoading","commentId":"M:AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading()","nameWithType":"PreloadedSceneHelper.FinishLoading()"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard","name":"Discard()","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_Discard","commentId":"M:AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard()","nameWithType":"PreloadedSceneHelper.Discard()"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.#ctor*","name":"PreloadedSceneHelper","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper__ctor_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.PreloadedSceneHelper","nameWithType":"PreloadedSceneHelper.PreloadedSceneHelper"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.scene*","name":"scene","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_scene_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.scene","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.scene","nameWithType":"PreloadedSceneHelper.scene"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded*","name":"isStillPreloaded","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_isStillPreloaded_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.isStillPreloaded","nameWithType":"PreloadedSceneHelper.isStillPreloaded"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks*","name":"hasRunCallbacks","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_hasRunCallbacks_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.hasRunCallbacks","nameWithType":"PreloadedSceneHelper.hasRunCallbacks"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading*","name":"FinishLoading","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_FinishLoading_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.FinishLoading","nameWithType":"PreloadedSceneHelper.FinishLoading"},{"uid":"AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard*","name":"Discard","href":"~/api/AdvancedSceneManager.Utility.PreloadedSceneHelper.yml#AdvancedSceneManager_Utility_PreloadedSceneHelper_Discard_","commentId":"Overload:AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard","isSpec":"True","fullName":"AdvancedSceneManager.Utility.PreloadedSceneHelper.Discard","nameWithType":"PreloadedSceneHelper.Discard"}],"api/AdvancedSceneManager.Utility.QueueUtility-1.yml":[{"uid":"AdvancedSceneManager.Utility.QueueUtility`1","name":"QueueUtility<T>","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml","commentId":"T:AdvancedSceneManager.Utility.QueueUtility`1","name.vb":"QueueUtility(Of T)","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T)","nameWithType":"QueueUtility<T>","nameWithType.vb":"QueueUtility(Of T)"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.isBusy","name":"isBusy","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_isBusy","commentId":"P:AdvancedSceneManager.Utility.QueueUtility`1.isBusy","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.isBusy","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).isBusy","nameWithType":"QueueUtility<T>.isBusy","nameWithType.vb":"QueueUtility(Of T).isBusy"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.queueEmpty","name":"queueEmpty","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_queueEmpty","commentId":"E:AdvancedSceneManager.Utility.QueueUtility`1.queueEmpty","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.queueEmpty","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).queueEmpty","nameWithType":"QueueUtility<T>.queueEmpty","nameWithType.vb":"QueueUtility(Of T).queueEmpty"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.queue","name":"queue","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_queue","commentId":"P:AdvancedSceneManager.Utility.QueueUtility`1.queue","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.queue","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).queue","nameWithType":"QueueUtility<T>.queue","nameWithType.vb":"QueueUtility(Of T).queue"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.running","name":"running","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_running","commentId":"P:AdvancedSceneManager.Utility.QueueUtility`1.running","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.running","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).running","nameWithType":"QueueUtility<T>.running","nameWithType.vb":"QueueUtility(Of T).running"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.IsQueued(`0)","name":"IsQueued(T)","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_IsQueued__0_","commentId":"M:AdvancedSceneManager.Utility.QueueUtility`1.IsQueued(`0)","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.IsQueued(T)","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).IsQueued(T)","nameWithType":"QueueUtility<T>.IsQueued(T)","nameWithType.vb":"QueueUtility(Of T).IsQueued(T)"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.IsRunning(`0)","name":"IsRunning(T)","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_IsRunning__0_","commentId":"M:AdvancedSceneManager.Utility.QueueUtility`1.IsRunning(`0)","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.IsRunning(T)","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).IsRunning(T)","nameWithType":"QueueUtility<T>.IsRunning(T)","nameWithType.vb":"QueueUtility(Of T).IsRunning(T)"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.StopAll","name":"StopAll()","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_StopAll","commentId":"M:AdvancedSceneManager.Utility.QueueUtility`1.StopAll","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.StopAll()","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).StopAll()","nameWithType":"QueueUtility<T>.StopAll()","nameWithType.vb":"QueueUtility(Of T).StopAll()"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.isBusy*","name":"isBusy","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_isBusy_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.isBusy","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.isBusy","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).isBusy","nameWithType":"QueueUtility<T>.isBusy","nameWithType.vb":"QueueUtility(Of T).isBusy"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.queue*","name":"queue","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_queue_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.queue","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.queue","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).queue","nameWithType":"QueueUtility<T>.queue","nameWithType.vb":"QueueUtility(Of T).queue"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.running*","name":"running","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_running_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.running","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.running","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).running","nameWithType":"QueueUtility<T>.running","nameWithType.vb":"QueueUtility(Of T).running"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.IsQueued*","name":"IsQueued","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_IsQueued_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.IsQueued","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.IsQueued","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).IsQueued","nameWithType":"QueueUtility<T>.IsQueued","nameWithType.vb":"QueueUtility(Of T).IsQueued"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.IsRunning*","name":"IsRunning","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_IsRunning_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.IsRunning","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.IsRunning","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).IsRunning","nameWithType":"QueueUtility<T>.IsRunning","nameWithType.vb":"QueueUtility(Of T).IsRunning"},{"uid":"AdvancedSceneManager.Utility.QueueUtility`1.StopAll*","name":"StopAll","href":"~/api/AdvancedSceneManager.Utility.QueueUtility-1.yml#AdvancedSceneManager_Utility_QueueUtility_1_StopAll_","commentId":"Overload:AdvancedSceneManager.Utility.QueueUtility`1.StopAll","isSpec":"True","fullName":"AdvancedSceneManager.Utility.QueueUtility<T>.StopAll","fullName.vb":"AdvancedSceneManager.Utility.QueueUtility(Of T).StopAll","nameWithType":"QueueUtility<T>.StopAll","nameWithType.vb":"QueueUtility(Of T).StopAll"}],"api/AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.yml":[{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode","name":"CallbackUtility.ShowMode","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.yml","commentId":"T:AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode","nameWithType":"CallbackUtility.ShowMode"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Time","name":"Time","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.yml#AdvancedSceneManager_Callbacks_CallbackUtility_ShowMode_Time","commentId":"F:AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Time","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Time","nameWithType":"CallbackUtility.ShowMode.Time"},{"uid":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Frames","name":"Frames","href":"~/api/AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.yml#AdvancedSceneManager_Callbacks_CallbackUtility_ShowMode_Frames","commentId":"F:AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Frames","fullName":"AdvancedSceneManager.Callbacks.CallbackUtility.ShowMode.Frames","nameWithType":"CallbackUtility.ShowMode.Frames"}],"api/AdvancedSceneManager.Core.SceneOperation.yml":[{"uid":"AdvancedSceneManager.Core.SceneOperation","name":"SceneOperation","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml","commentId":"T:AdvancedSceneManager.Core.SceneOperation","fullName":"AdvancedSceneManager.Core.SceneOperation","nameWithType":"SceneOperation"},{"uid":"AdvancedSceneManager.Core.SceneOperation.done","name":"done","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_done","commentId":"P:AdvancedSceneManager.Core.SceneOperation.done","fullName":"AdvancedSceneManager.Core.SceneOperation.done","nameWithType":"SceneOperation.done"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Add(AdvancedSceneManager.Core.SceneManagerBase,System.Boolean)","name":"Add(SceneManagerBase, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Add_AdvancedSceneManager_Core_SceneManagerBase_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Add(AdvancedSceneManager.Core.SceneManagerBase,System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.Add(AdvancedSceneManager.Core.SceneManagerBase, System.Boolean)","nameWithType":"SceneOperation.Add(SceneManagerBase, Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Add``1(AdvancedSceneManager.Core.SceneManagerBase,System.Boolean)","name":"Add<ReturnValue>(SceneManagerBase, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Add__1_AdvancedSceneManager_Core_SceneManagerBase_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Add``1(AdvancedSceneManager.Core.SceneManagerBase,System.Boolean)","name.vb":"Add(Of ReturnValue)(SceneManagerBase, Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.Add<ReturnValue>(AdvancedSceneManager.Core.SceneManagerBase, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Add(Of ReturnValue)(AdvancedSceneManager.Core.SceneManagerBase, System.Boolean)","nameWithType":"SceneOperation.Add<ReturnValue>(SceneManagerBase, Boolean)","nameWithType.vb":"SceneOperation.Add(Of ReturnValue)(SceneManagerBase, Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Add``1(AdvancedSceneManager.Core.SceneManagerBase,System.Func{AdvancedSceneManager.Core.SceneOperation,``0},System.Boolean)","name":"Add<ReturnValue>(SceneManagerBase, Func<SceneOperation, ReturnValue>, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Add__1_AdvancedSceneManager_Core_SceneManagerBase_System_Func_AdvancedSceneManager_Core_SceneOperation___0__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Add``1(AdvancedSceneManager.Core.SceneManagerBase,System.Func{AdvancedSceneManager.Core.SceneOperation,``0},System.Boolean)","name.vb":"Add(Of ReturnValue)(SceneManagerBase, Func(Of SceneOperation, ReturnValue), Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.Add<ReturnValue>(AdvancedSceneManager.Core.SceneManagerBase, System.Func<AdvancedSceneManager.Core.SceneOperation, ReturnValue>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Add(Of ReturnValue)(AdvancedSceneManager.Core.SceneManagerBase, System.Func(Of AdvancedSceneManager.Core.SceneOperation, ReturnValue), System.Boolean)","nameWithType":"SceneOperation.Add<ReturnValue>(SceneManagerBase, Func<SceneOperation, ReturnValue>, Boolean)","nameWithType.vb":"SceneOperation.Add(Of ReturnValue)(SceneManagerBase, Func(Of SceneOperation, ReturnValue), Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnTurn(System.Action)","name":"IQueueable.OnTurn(Action)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AdvancedSceneManager_Utility_IQueueable_OnTurn_System_Action_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnTurn(System.Action)","name.vb":"AdvancedSceneManager.Utility.IQueueable.OnTurn(Action)","fullName":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnTurn(System.Action)","nameWithType":"SceneOperation.IQueueable.OnTurn(Action)","nameWithType.vb":"SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnTurn(Action)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnCancel","name":"IQueueable.OnCancel()","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AdvancedSceneManager_Utility_IQueueable_OnCancel","commentId":"M:AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnCancel","name.vb":"AdvancedSceneManager.Utility.IQueueable.OnCancel()","fullName":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnCancel()","nameWithType":"SceneOperation.IQueueable.OnCancel()","nameWithType.vb":"SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnCancel()"},{"uid":"AdvancedSceneManager.Core.SceneOperation.friendlyText","name":"friendlyText","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_friendlyText","commentId":"P:AdvancedSceneManager.Core.SceneOperation.friendlyText","fullName":"AdvancedSceneManager.Core.SceneOperation.friendlyText","nameWithType":"SceneOperation.friendlyText"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithFriendlyText(System.String)","name":"WithFriendlyText(String)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithFriendlyText_System_String_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithFriendlyText(System.String)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithFriendlyText(System.String)","nameWithType":"SceneOperation.WithFriendlyText(String)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.open","name":"open","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_open","commentId":"P:AdvancedSceneManager.Core.SceneOperation.open","fullName":"AdvancedSceneManager.Core.SceneOperation.open","nameWithType":"SceneOperation.open"},{"uid":"AdvancedSceneManager.Core.SceneOperation.close","name":"close","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_close","commentId":"P:AdvancedSceneManager.Core.SceneOperation.close","fullName":"AdvancedSceneManager.Core.SceneOperation.close","nameWithType":"SceneOperation.close"},{"uid":"AdvancedSceneManager.Core.SceneOperation.reopen","name":"reopen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_reopen","commentId":"P:AdvancedSceneManager.Core.SceneOperation.reopen","fullName":"AdvancedSceneManager.Core.SceneOperation.reopen","nameWithType":"SceneOperation.reopen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.customActions","name":"customActions","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_customActions","commentId":"P:AdvancedSceneManager.Core.SceneOperation.customActions","fullName":"AdvancedSceneManager.Core.SceneOperation.customActions","nameWithType":"SceneOperation.customActions"},{"uid":"AdvancedSceneManager.Core.SceneOperation.callbacks","name":"callbacks","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_callbacks","commentId":"P:AdvancedSceneManager.Core.SceneOperation.callbacks","fullName":"AdvancedSceneManager.Core.SceneOperation.callbacks","nameWithType":"SceneOperation.callbacks"},{"uid":"AdvancedSceneManager.Core.SceneOperation.collection","name":"collection","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_collection","commentId":"P:AdvancedSceneManager.Core.SceneOperation.collection","fullName":"AdvancedSceneManager.Core.SceneOperation.collection","nameWithType":"SceneOperation.collection"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingScreen","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingScreen","commentId":"P:AdvancedSceneManager.Core.SceneOperation.loadingScreen","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingScreen","nameWithType":"SceneOperation.loadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.useLoadingScreen","name":"useLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_useLoadingScreen","commentId":"P:AdvancedSceneManager.Core.SceneOperation.useLoadingScreen","fullName":"AdvancedSceneManager.Core.SceneOperation.useLoadingScreen","nameWithType":"SceneOperation.useLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets","name":"clearUnusedAssets","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_clearUnusedAssets","commentId":"P:AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets","fullName":"AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets","nameWithType":"SceneOperation.clearUnusedAssets"},{"uid":"AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks","name":"doCollectionCallbacks","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_doCollectionCallbacks","commentId":"P:AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks","fullName":"AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks","nameWithType":"SceneOperation.doCollectionCallbacks"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback","name":"loadingScreenCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingScreenCallback","commentId":"P:AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback","nameWithType":"SceneOperation.loadingScreenCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingPriority","name":"loadingPriority","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingPriority","commentId":"P:AdvancedSceneManager.Core.SceneOperation.loadingPriority","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingPriority","nameWithType":"SceneOperation.loadingPriority"},{"uid":"AdvancedSceneManager.Core.SceneOperation.closeBehavior","name":"closeBehavior","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_closeBehavior","commentId":"P:AdvancedSceneManager.Core.SceneOperation.closeBehavior","fullName":"AdvancedSceneManager.Core.SceneOperation.closeBehavior","nameWithType":"SceneOperation.closeBehavior"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Open(AdvancedSceneManager.Models.Scene[])","name":"Open(Scene[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Open_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Open(AdvancedSceneManager.Models.Scene[])","name.vb":"Open(Scene())","fullName":"AdvancedSceneManager.Core.SceneOperation.Open(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Open(AdvancedSceneManager.Models.Scene())","nameWithType":"SceneOperation.Open(Scene[])","nameWithType.vb":"SceneOperation.Open(Scene())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Open(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.Boolean)","name":"Open(IEnumerable<Scene>, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Open_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Models_Scene__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Open(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene},System.Boolean)","name.vb":"Open(IEnumerable(Of Scene), Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.Open(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Models.Scene>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Open(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Models.Scene), System.Boolean)","nameWithType":"SceneOperation.Open(IEnumerable<Scene>, Boolean)","nameWithType.vb":"SceneOperation.Open(IEnumerable(Of Scene), Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Close(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Close_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Close(OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation.Close(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Close(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation.Close(OpenSceneInfo[])","nameWithType.vb":"SceneOperation.Close(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Close(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},System.Boolean)","name":"Close(IEnumerable<OpenSceneInfo>, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Close_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Close(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo},System.Boolean)","name.vb":"Close(IEnumerable(Of OpenSceneInfo), Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.Close(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>, System.Boolean)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Close(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo), System.Boolean)","nameWithType":"SceneOperation.Close(IEnumerable<OpenSceneInfo>, Boolean)","nameWithType.vb":"SceneOperation.Close(IEnumerable(Of OpenSceneInfo), Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Close(System.Boolean,AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Close(Boolean, OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Close_System_Boolean_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Close(System.Boolean,AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Close(Boolean, OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation.Close(System.Boolean, AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Close(System.Boolean, AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation.Close(Boolean, OpenSceneInfo[])","nameWithType.vb":"SceneOperation.Close(Boolean, OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","name":"Reopen(OpenSceneInfo[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Reopen_AdvancedSceneManager_Core_OpenSceneInfo___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","name.vb":"Reopen(OpenSceneInfo())","fullName":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Core.OpenSceneInfo[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Core.OpenSceneInfo())","nameWithType":"SceneOperation.Reopen(OpenSceneInfo[])","nameWithType.vb":"SceneOperation.Reopen(OpenSceneInfo())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo})","name":"Reopen(IEnumerable<OpenSceneInfo>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Reopen_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Core_OpenSceneInfo__","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Core.OpenSceneInfo})","name.vb":"Reopen(IEnumerable(Of OpenSceneInfo))","fullName":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Core.OpenSceneInfo>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Core.OpenSceneInfo))","nameWithType":"SceneOperation.Reopen(IEnumerable<OpenSceneInfo>)","nameWithType.vb":"SceneOperation.Reopen(IEnumerable(Of OpenSceneInfo))"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Models.Scene[])","name":"Reopen(Scene[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Reopen_AdvancedSceneManager_Models_Scene___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Models.Scene[])","name.vb":"Reopen(Scene())","fullName":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Models.Scene[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Reopen(AdvancedSceneManager.Models.Scene())","nameWithType":"SceneOperation.Reopen(Scene[])","nameWithType.vb":"SceneOperation.Reopen(Scene())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene})","name":"Reopen(IEnumerable<Scene>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Reopen_System_Collections_Generic_IEnumerable_AdvancedSceneManager_Models_Scene__","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable{AdvancedSceneManager.Models.Scene})","name.vb":"Reopen(IEnumerable(Of Scene))","fullName":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable<AdvancedSceneManager.Models.Scene>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.Reopen(System.Collections.Generic.IEnumerable(Of AdvancedSceneManager.Models.Scene))","nameWithType":"SceneOperation.Reopen(IEnumerable<Scene>)","nameWithType.vb":"SceneOperation.Reopen(IEnumerable(Of Scene))"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","name":"WithAction(SceneAction[])","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithAction_AdvancedSceneManager_Core_Actions_SceneAction___","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","name.vb":"WithAction(SceneAction())","fullName":"AdvancedSceneManager.Core.SceneOperation.WithAction(AdvancedSceneManager.Core.Actions.SceneAction[])","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.WithAction(AdvancedSceneManager.Core.Actions.SceneAction())","nameWithType":"SceneOperation.WithAction(SceneAction[])","nameWithType.vb":"SceneOperation.WithAction(SceneAction())"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithCallback(AdvancedSceneManager.Core.Callback)","name":"WithCallback(Callback)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithCallback_AdvancedSceneManager_Core_Callback_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithCallback(AdvancedSceneManager.Core.Callback)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithCallback(AdvancedSceneManager.Core.Callback)","nameWithType":"SceneOperation.WithCallback(Callback)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithCollection(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","name":"WithCollection(SceneCollection, Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithCollection_AdvancedSceneManager_Models_SceneCollection_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithCollection(AdvancedSceneManager.Models.SceneCollection,System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithCollection(AdvancedSceneManager.Models.SceneCollection, System.Boolean)","nameWithType":"SceneOperation.WithCollection(SceneCollection, Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(System.Boolean)","name":"WithLoadingScreen(Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingScreen_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(System.Boolean)","nameWithType":"SceneOperation.WithLoadingScreen(Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","name":"WithLoadingScreen(Scene)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingScreen_AdvancedSceneManager_Models_Scene_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen(AdvancedSceneManager.Models.Scene)","nameWithType":"SceneOperation.WithLoadingScreen(Scene)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets(System.Boolean)","name":"WithClearUnusedAssets(Boolean)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithClearUnusedAssets_System_Boolean_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets(System.Boolean)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets(System.Boolean)","nameWithType":"SceneOperation.WithClearUnusedAssets(Boolean)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback(System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name":"WithLoadingScreenCallback(Action<LoadingScreen>)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingScreenCallback_System_Action_AdvancedSceneManager_Callbacks_LoadingScreen__","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback(System.Action{AdvancedSceneManager.Callbacks.LoadingScreen})","name.vb":"WithLoadingScreenCallback(Action(Of LoadingScreen))","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback(System.Action<AdvancedSceneManager.Callbacks.LoadingScreen>)","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback(System.Action(Of AdvancedSceneManager.Callbacks.LoadingScreen))","nameWithType":"SceneOperation.WithLoadingScreenCallback(Action<LoadingScreen>)","nameWithType.vb":"SceneOperation.WithLoadingScreenCallback(Action(Of LoadingScreen))"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority(UnityEngine.ThreadPriority)","name":"WithLoadingPriority(ThreadPriority)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingPriority_UnityEngine_ThreadPriority_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority(UnityEngine.ThreadPriority)","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority(UnityEngine.ThreadPriority)","nameWithType":"SceneOperation.WithLoadingPriority(ThreadPriority)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","name":"AsPersistent(SceneCloseBehavior)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AsPersistent_AdvancedSceneManager_Models_SceneCloseBehavior_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","fullName":"AdvancedSceneManager.Core.SceneOperation.AsPersistent(AdvancedSceneManager.Models.SceneCloseBehavior)","nameWithType":"SceneOperation.AsPersistent(SceneCloseBehavior)"},{"uid":"AdvancedSceneManager.Core.SceneOperation._extCallbacks","name":"_extCallbacks","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation__extCallbacks","commentId":"F:AdvancedSceneManager.Core.SceneOperation._extCallbacks","fullName":"AdvancedSceneManager.Core.SceneOperation._extCallbacks","nameWithType":"SceneOperation._extCallbacks"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AddCallback(AdvancedSceneManager.Core.Callback)","name":"AddCallback(Callback)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AddCallback_AdvancedSceneManager_Core_Callback_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.AddCallback(AdvancedSceneManager.Core.Callback)","fullName":"AdvancedSceneManager.Core.SceneOperation.AddCallback(AdvancedSceneManager.Core.Callback)","nameWithType":"SceneOperation.AddCallback(Callback)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.RemoveCallback(AdvancedSceneManager.Core.Callback)","name":"RemoveCallback(Callback)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_RemoveCallback_AdvancedSceneManager_Core_Callback_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.RemoveCallback(AdvancedSceneManager.Core.Callback)","fullName":"AdvancedSceneManager.Core.SceneOperation.RemoveCallback(AdvancedSceneManager.Core.Callback)","nameWithType":"SceneOperation.RemoveCallback(Callback)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.keepWaiting","name":"keepWaiting","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_keepWaiting","commentId":"P:AdvancedSceneManager.Core.SceneOperation.keepWaiting","fullName":"AdvancedSceneManager.Core.SceneOperation.keepWaiting","nameWithType":"SceneOperation.keepWaiting"},{"uid":"AdvancedSceneManager.Core.SceneOperation.phase","name":"phase","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_phase","commentId":"P:AdvancedSceneManager.Core.SceneOperation.phase","fullName":"AdvancedSceneManager.Core.SceneOperation.phase","nameWithType":"SceneOperation.phase"},{"uid":"AdvancedSceneManager.Core.SceneOperation.sceneManager","name":"sceneManager","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_sceneManager","commentId":"P:AdvancedSceneManager.Core.SceneOperation.sceneManager","fullName":"AdvancedSceneManager.Core.SceneOperation.sceneManager","nameWithType":"SceneOperation.sceneManager"},{"uid":"AdvancedSceneManager.Core.SceneOperation.current","name":"current","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_current","commentId":"P:AdvancedSceneManager.Core.SceneOperation.current","fullName":"AdvancedSceneManager.Core.SceneOperation.current","nameWithType":"SceneOperation.current"},{"uid":"AdvancedSceneManager.Core.SceneOperation.cancelled","name":"cancelled","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_cancelled","commentId":"P:AdvancedSceneManager.Core.SceneOperation.cancelled","fullName":"AdvancedSceneManager.Core.SceneOperation.cancelled","nameWithType":"SceneOperation.cancelled"},{"uid":"AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen","name":"openedLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_openedLoadingScreen","commentId":"P:AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen","fullName":"AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen","nameWithType":"SceneOperation.openedLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.actions","name":"actions","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_actions","commentId":"P:AdvancedSceneManager.Core.SceneOperation.actions","fullName":"AdvancedSceneManager.Core.SceneOperation.actions","nameWithType":"SceneOperation.actions"},{"uid":"AdvancedSceneManager.Core.SceneOperation.totalProgress","name":"totalProgress","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_totalProgress","commentId":"P:AdvancedSceneManager.Core.SceneOperation.totalProgress","fullName":"AdvancedSceneManager.Core.SceneOperation.totalProgress","nameWithType":"SceneOperation.totalProgress"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Cancel(System.Action)","name":"Cancel(Action)","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Cancel_System_Action_","commentId":"M:AdvancedSceneManager.Core.SceneOperation.Cancel(System.Action)","fullName":"AdvancedSceneManager.Core.SceneOperation.Cancel(System.Action)","nameWithType":"SceneOperation.Cancel(Action)"},{"uid":"AdvancedSceneManager.Core.SceneOperation.isDone","name":"isDone","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_isDone","commentId":"F:AdvancedSceneManager.Core.SceneOperation.isDone","fullName":"AdvancedSceneManager.Core.SceneOperation.isDone","nameWithType":"SceneOperation.isDone"},{"uid":"AdvancedSceneManager.Core.SceneOperation.FindActions``1","name":"FindActions<T>()","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_FindActions__1","commentId":"M:AdvancedSceneManager.Core.SceneOperation.FindActions``1","name.vb":"FindActions(Of T)()","fullName":"AdvancedSceneManager.Core.SceneOperation.FindActions<T>()","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.FindActions(Of T)()","nameWithType":"SceneOperation.FindActions<T>()","nameWithType.vb":"SceneOperation.FindActions(Of T)()"},{"uid":"AdvancedSceneManager.Core.SceneOperation.FindLastAction``1","name":"FindLastAction<T>()","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_FindLastAction__1","commentId":"M:AdvancedSceneManager.Core.SceneOperation.FindLastAction``1","name.vb":"FindLastAction(Of T)()","fullName":"AdvancedSceneManager.Core.SceneOperation.FindLastAction<T>()","fullName.vb":"AdvancedSceneManager.Core.SceneOperation.FindLastAction(Of T)()","nameWithType":"SceneOperation.FindLastAction<T>()","nameWithType.vb":"SceneOperation.FindLastAction(Of T)()"},{"uid":"AdvancedSceneManager.Core.SceneOperation.openedScenes","name":"openedScenes","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_openedScenes","commentId":"P:AdvancedSceneManager.Core.SceneOperation.openedScenes","fullName":"AdvancedSceneManager.Core.SceneOperation.openedScenes","nameWithType":"SceneOperation.openedScenes"},{"uid":"AdvancedSceneManager.Core.SceneOperation.done*","name":"done","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_done_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.done","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.done","nameWithType":"SceneOperation.done"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Add*","name":"Add","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Add_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.Add","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.Add","nameWithType":"SceneOperation.Add"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnTurn*","name":"IQueueable.OnTurn","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AdvancedSceneManager_Utility_IQueueable_OnTurn_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnTurn","isSpec":"True","name.vb":"AdvancedSceneManager.Utility.IQueueable.OnTurn","fullName":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnTurn","nameWithType":"SceneOperation.IQueueable.OnTurn","nameWithType.vb":"SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnTurn"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnCancel*","name":"IQueueable.OnCancel","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AdvancedSceneManager_Utility_IQueueable_OnCancel_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager#Utility#IQueueable#OnCancel","isSpec":"True","name.vb":"AdvancedSceneManager.Utility.IQueueable.OnCancel","fullName":"AdvancedSceneManager.Core.SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnCancel","nameWithType":"SceneOperation.IQueueable.OnCancel","nameWithType.vb":"SceneOperation.AdvancedSceneManager.Utility.IQueueable.OnCancel"},{"uid":"AdvancedSceneManager.Core.SceneOperation.friendlyText*","name":"friendlyText","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_friendlyText_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.friendlyText","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.friendlyText","nameWithType":"SceneOperation.friendlyText"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithFriendlyText*","name":"WithFriendlyText","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithFriendlyText_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithFriendlyText","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithFriendlyText","nameWithType":"SceneOperation.WithFriendlyText"},{"uid":"AdvancedSceneManager.Core.SceneOperation.open*","name":"open","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_open_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.open","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.open","nameWithType":"SceneOperation.open"},{"uid":"AdvancedSceneManager.Core.SceneOperation.close*","name":"close","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_close_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.close","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.close","nameWithType":"SceneOperation.close"},{"uid":"AdvancedSceneManager.Core.SceneOperation.reopen*","name":"reopen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_reopen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.reopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.reopen","nameWithType":"SceneOperation.reopen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.customActions*","name":"customActions","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_customActions_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.customActions","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.customActions","nameWithType":"SceneOperation.customActions"},{"uid":"AdvancedSceneManager.Core.SceneOperation.callbacks*","name":"callbacks","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_callbacks_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.callbacks","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.callbacks","nameWithType":"SceneOperation.callbacks"},{"uid":"AdvancedSceneManager.Core.SceneOperation.collection*","name":"collection","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_collection_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.collection","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.collection","nameWithType":"SceneOperation.collection"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingScreen*","name":"loadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.loadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingScreen","nameWithType":"SceneOperation.loadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.useLoadingScreen*","name":"useLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_useLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.useLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.useLoadingScreen","nameWithType":"SceneOperation.useLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets*","name":"clearUnusedAssets","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_clearUnusedAssets_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.clearUnusedAssets","nameWithType":"SceneOperation.clearUnusedAssets"},{"uid":"AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks*","name":"doCollectionCallbacks","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_doCollectionCallbacks_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.doCollectionCallbacks","nameWithType":"SceneOperation.doCollectionCallbacks"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback*","name":"loadingScreenCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingScreenCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingScreenCallback","nameWithType":"SceneOperation.loadingScreenCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.loadingPriority*","name":"loadingPriority","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_loadingPriority_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.loadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.loadingPriority","nameWithType":"SceneOperation.loadingPriority"},{"uid":"AdvancedSceneManager.Core.SceneOperation.closeBehavior*","name":"closeBehavior","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_closeBehavior_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.closeBehavior","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.closeBehavior","nameWithType":"SceneOperation.closeBehavior"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Open_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.Open","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.Open","nameWithType":"SceneOperation.Open"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Close_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.Close","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.Close","nameWithType":"SceneOperation.Close"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Reopen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.Reopen","nameWithType":"SceneOperation.Reopen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithAction*","name":"WithAction","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithAction_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithAction","nameWithType":"SceneOperation.WithAction"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithCallback*","name":"WithCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithCallback","nameWithType":"SceneOperation.WithCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithCollection*","name":"WithCollection","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithCollection_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithCollection","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithCollection","nameWithType":"SceneOperation.WithCollection"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen*","name":"WithLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreen","nameWithType":"SceneOperation.WithLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets*","name":"WithClearUnusedAssets","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithClearUnusedAssets_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithClearUnusedAssets","nameWithType":"SceneOperation.WithClearUnusedAssets"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback*","name":"WithLoadingScreenCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingScreenCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingScreenCallback","nameWithType":"SceneOperation.WithLoadingScreenCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority*","name":"WithLoadingPriority","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_WithLoadingPriority_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.WithLoadingPriority","nameWithType":"SceneOperation.WithLoadingPriority"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AsPersistent*","name":"AsPersistent","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AsPersistent_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.AsPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.AsPersistent","nameWithType":"SceneOperation.AsPersistent"},{"uid":"AdvancedSceneManager.Core.SceneOperation.AddCallback*","name":"AddCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_AddCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.AddCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.AddCallback","nameWithType":"SceneOperation.AddCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.RemoveCallback*","name":"RemoveCallback","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_RemoveCallback_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.RemoveCallback","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.RemoveCallback","nameWithType":"SceneOperation.RemoveCallback"},{"uid":"AdvancedSceneManager.Core.SceneOperation.keepWaiting*","name":"keepWaiting","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_keepWaiting_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.keepWaiting","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.keepWaiting","nameWithType":"SceneOperation.keepWaiting"},{"uid":"AdvancedSceneManager.Core.SceneOperation.phase*","name":"phase","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_phase_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.phase","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.phase","nameWithType":"SceneOperation.phase"},{"uid":"AdvancedSceneManager.Core.SceneOperation.sceneManager*","name":"sceneManager","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_sceneManager_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.sceneManager","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.sceneManager","nameWithType":"SceneOperation.sceneManager"},{"uid":"AdvancedSceneManager.Core.SceneOperation.current*","name":"current","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_current_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.current","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.current","nameWithType":"SceneOperation.current"},{"uid":"AdvancedSceneManager.Core.SceneOperation.cancelled*","name":"cancelled","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_cancelled_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.cancelled","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.cancelled","nameWithType":"SceneOperation.cancelled"},{"uid":"AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen*","name":"openedLoadingScreen","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_openedLoadingScreen_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.openedLoadingScreen","nameWithType":"SceneOperation.openedLoadingScreen"},{"uid":"AdvancedSceneManager.Core.SceneOperation.actions*","name":"actions","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_actions_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.actions","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.actions","nameWithType":"SceneOperation.actions"},{"uid":"AdvancedSceneManager.Core.SceneOperation.totalProgress*","name":"totalProgress","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_totalProgress_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.totalProgress","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.totalProgress","nameWithType":"SceneOperation.totalProgress"},{"uid":"AdvancedSceneManager.Core.SceneOperation.Cancel*","name":"Cancel","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_Cancel_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.Cancel","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.Cancel","nameWithType":"SceneOperation.Cancel"},{"uid":"AdvancedSceneManager.Core.SceneOperation.FindActions*","name":"FindActions","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_FindActions_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.FindActions","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.FindActions","nameWithType":"SceneOperation.FindActions"},{"uid":"AdvancedSceneManager.Core.SceneOperation.FindLastAction*","name":"FindLastAction","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_FindLastAction_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.FindLastAction","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.FindLastAction","nameWithType":"SceneOperation.FindLastAction"},{"uid":"AdvancedSceneManager.Core.SceneOperation.openedScenes*","name":"openedScenes","href":"~/api/AdvancedSceneManager.Core.SceneOperation.yml#AdvancedSceneManager_Core_SceneOperation_openedScenes_","commentId":"Overload:AdvancedSceneManager.Core.SceneOperation.openedScenes","isSpec":"True","fullName":"AdvancedSceneManager.Core.SceneOperation.openedScenes","nameWithType":"SceneOperation.openedScenes"}],"api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml":[{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen","name":"IconBounceLoadingScreen","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml","commentId":"T:AdvancedSceneManager.Defaults.IconBounceLoadingScreen","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen","nameWithType":"IconBounceLoadingScreen"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartSize","name":"IconStartSize","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_IconStartSize","commentId":"F:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartSize","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartSize","nameWithType":"IconBounceLoadingScreen.IconStartSize"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartRotationZ","name":"IconStartRotationZ","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_IconStartRotationZ","commentId":"F:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartRotationZ","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconStartRotationZ","nameWithType":"IconBounceLoadingScreen.IconStartRotationZ"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.duration","name":"duration","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_duration","commentId":"F:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.duration","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.duration","nameWithType":"IconBounceLoadingScreen.duration"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconTransform","name":"IconTransform","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_IconTransform","commentId":"F:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconTransform","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.IconTransform","nameWithType":"IconBounceLoadingScreen.IconTransform"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.BackgroundTransform","name":"BackgroundTransform","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_BackgroundTransform","commentId":"F:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.BackgroundTransform","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.BackgroundTransform","nameWithType":"IconBounceLoadingScreen.BackgroundTransform"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","name":"OnOpen(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_OnOpen_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"IconBounceLoadingScreen.OnOpen(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","name":"OnClose(SceneOperation)","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_OnClose_AdvancedSceneManager_Core_SceneOperation_","commentId":"M:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose(AdvancedSceneManager.Core.SceneOperation)","nameWithType":"IconBounceLoadingScreen.OnClose(SceneOperation)"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen*","name":"OnOpen","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_OnOpen_","commentId":"Overload:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnOpen","nameWithType":"IconBounceLoadingScreen.OnOpen"},{"uid":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Defaults.IconBounceLoadingScreen.yml#AdvancedSceneManager_Defaults_IconBounceLoadingScreen_OnClose_","commentId":"Overload:AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Defaults.IconBounceLoadingScreen.OnClose","nameWithType":"IconBounceLoadingScreen.OnClose"}],"api/AdvancedSceneManager.Defaults.Quotes.Quote.yml":[{"uid":"AdvancedSceneManager.Defaults.Quotes.Quote","name":"Quotes.Quote","href":"~/api/AdvancedSceneManager.Defaults.Quotes.Quote.yml","commentId":"T:AdvancedSceneManager.Defaults.Quotes.Quote","fullName":"AdvancedSceneManager.Defaults.Quotes.Quote","nameWithType":"Quotes.Quote"},{"uid":"AdvancedSceneManager.Defaults.Quotes.Quote.name","name":"name","href":"~/api/AdvancedSceneManager.Defaults.Quotes.Quote.yml#AdvancedSceneManager_Defaults_Quotes_Quote_name","commentId":"F:AdvancedSceneManager.Defaults.Quotes.Quote.name","fullName":"AdvancedSceneManager.Defaults.Quotes.Quote.name","nameWithType":"Quotes.Quote.name"},{"uid":"AdvancedSceneManager.Defaults.Quotes.Quote.quote","name":"quote","href":"~/api/AdvancedSceneManager.Defaults.Quotes.Quote.yml#AdvancedSceneManager_Defaults_Quotes_Quote_quote","commentId":"F:AdvancedSceneManager.Defaults.Quotes.Quote.quote","fullName":"AdvancedSceneManager.Defaults.Quotes.Quote.quote","nameWithType":"Quotes.Quote.quote"}],"api/AdvancedSceneManager.Editor.GenericPopup.yml":[{"uid":"AdvancedSceneManager.Editor.GenericPopup","name":"GenericPopup","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml","commentId":"T:AdvancedSceneManager.Editor.GenericPopup","fullName":"AdvancedSceneManager.Editor.GenericPopup","nameWithType":"GenericPopup"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_path","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.path","fullName":"AdvancedSceneManager.Editor.GenericPopup.path","nameWithType":"GenericPopup.path"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Separator","name":"Separator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_Separator","commentId":"P:AdvancedSceneManager.Editor.GenericPopup.Separator","fullName":"AdvancedSceneManager.Editor.GenericPopup.Separator","nameWithType":"GenericPopup.Separator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Refresh(AdvancedSceneManager.Editor.GenericPopup.Item[])","name":"Refresh(GenericPopup.Item[])","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_Refresh_AdvancedSceneManager_Editor_GenericPopup_Item___","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.Refresh(AdvancedSceneManager.Editor.GenericPopup.Item[])","name.vb":"Refresh(GenericPopup.Item())","fullName":"AdvancedSceneManager.Editor.GenericPopup.Refresh(AdvancedSceneManager.Editor.GenericPopup.Item[])","fullName.vb":"AdvancedSceneManager.Editor.GenericPopup.Refresh(AdvancedSceneManager.Editor.GenericPopup.Item())","nameWithType":"GenericPopup.Refresh(GenericPopup.Item[])","nameWithType.vb":"GenericPopup.Refresh(GenericPopup.Item())"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.OnReopen(AdvancedSceneManager.Editor.GenericPopup)","name":"OnReopen(GenericPopup)","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_OnReopen_AdvancedSceneManager_Editor_GenericPopup_","commentId":"M:AdvancedSceneManager.Editor.GenericPopup.OnReopen(AdvancedSceneManager.Editor.GenericPopup)","fullName":"AdvancedSceneManager.Editor.GenericPopup.OnReopen(AdvancedSceneManager.Editor.GenericPopup)","nameWithType":"GenericPopup.OnReopen(GenericPopup)"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_path_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.path","nameWithType":"GenericPopup.path"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Separator*","name":"Separator","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_Separator_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Separator","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Separator","nameWithType":"GenericPopup.Separator"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.Refresh*","name":"Refresh","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_Refresh_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.Refresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.Refresh","nameWithType":"GenericPopup.Refresh"},{"uid":"AdvancedSceneManager.Editor.GenericPopup.OnReopen*","name":"OnReopen","href":"~/api/AdvancedSceneManager.Editor.GenericPopup.yml#AdvancedSceneManager_Editor_GenericPopup_OnReopen_","commentId":"Overload:AdvancedSceneManager.Editor.GenericPopup.OnReopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.GenericPopup.OnReopen","nameWithType":"GenericPopup.OnReopen"}],"api/AdvancedSceneManager.Editor.Popup-1.yml":[{"uid":"AdvancedSceneManager.Editor.Popup`1","name":"Popup<T>","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml","commentId":"T:AdvancedSceneManager.Editor.Popup`1","name.vb":"Popup(Of T)","fullName":"AdvancedSceneManager.Editor.Popup<T>","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T)","nameWithType":"Popup<T>","nameWithType.vb":"Popup(Of T)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Reopen","name":"Reopen()","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Reopen","commentId":"M:AdvancedSceneManager.Editor.Popup`1.Reopen","fullName":"AdvancedSceneManager.Editor.Popup<T>.Reopen()","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Reopen()","nameWithType":"Popup<T>.Reopen()","nameWithType.vb":"Popup(Of T).Reopen()"},{"uid":"AdvancedSceneManager.Editor.Popup`1.OnReopen(`0)","name":"OnReopen(T)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_OnReopen__0_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.OnReopen(`0)","fullName":"AdvancedSceneManager.Editor.Popup<T>.OnReopen(T)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).OnReopen(T)","nameWithType":"Popup<T>.OnReopen(T)","nameWithType.vb":"Popup(Of T).OnReopen(T)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Open(UnityEngine.UIElements.VisualElement,AdvancedSceneManager.Editor.IUIToolkitEditor,System.Boolean,UnityEngine.Vector2,System.Boolean,System.Boolean)","name":"Open(VisualElement, IUIToolkitEditor, Boolean, Vector2, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Open_UnityEngine_UIElements_VisualElement_AdvancedSceneManager_Editor_IUIToolkitEditor_System_Boolean_UnityEngine_Vector2_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.Open(UnityEngine.UIElements.VisualElement,AdvancedSceneManager.Editor.IUIToolkitEditor,System.Boolean,UnityEngine.Vector2,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Editor.Popup<T>.Open(UnityEngine.UIElements.VisualElement, AdvancedSceneManager.Editor.IUIToolkitEditor, System.Boolean, UnityEngine.Vector2, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Open(UnityEngine.UIElements.VisualElement, AdvancedSceneManager.Editor.IUIToolkitEditor, System.Boolean, UnityEngine.Vector2, System.Boolean, System.Boolean)","nameWithType":"Popup<T>.Open(VisualElement, IUIToolkitEditor, Boolean, Vector2, Boolean, Boolean)","nameWithType.vb":"Popup(Of T).Open(VisualElement, IUIToolkitEditor, Boolean, Vector2, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.CloseWithoutAnimation(System.Boolean)","name":"CloseWithoutAnimation(Boolean)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_CloseWithoutAnimation_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.CloseWithoutAnimation(System.Boolean)","fullName":"AdvancedSceneManager.Editor.Popup<T>.CloseWithoutAnimation(System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).CloseWithoutAnimation(System.Boolean)","nameWithType":"Popup<T>.CloseWithoutAnimation(Boolean)","nameWithType.vb":"Popup(Of T).CloseWithoutAnimation(Boolean)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Close","name":"Close()","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Close","commentId":"M:AdvancedSceneManager.Editor.Popup`1.Close","fullName":"AdvancedSceneManager.Editor.Popup<T>.Close()","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Close()","nameWithType":"Popup<T>.Close()","nameWithType.vb":"Popup(Of T).Close()"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Close(System.Action)","name":"Close(Action)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Close_System_Action_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.Close(System.Action)","fullName":"AdvancedSceneManager.Editor.Popup<T>.Close(System.Action)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Close(System.Action)","nameWithType":"Popup<T>.Close(Action)","nameWithType.vb":"Popup(Of T).Close(Action)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.OnClose","name":"OnClose()","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_OnClose","commentId":"M:AdvancedSceneManager.Editor.Popup`1.OnClose","fullName":"AdvancedSceneManager.Editor.Popup<T>.OnClose()","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).OnClose()","nameWithType":"Popup<T>.OnClose()","nameWithType.vb":"Popup(Of T).OnClose()"},{"uid":"AdvancedSceneManager.Editor.Popup`1.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_path","commentId":"P:AdvancedSceneManager.Editor.Popup`1.path","fullName":"AdvancedSceneManager.Editor.Popup<T>.path","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).path","nameWithType":"Popup<T>.path","nameWithType.vb":"Popup(Of T).path"},{"uid":"AdvancedSceneManager.Editor.Popup`1.overlay","name":"overlay","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_overlay","commentId":"F:AdvancedSceneManager.Editor.Popup`1.overlay","fullName":"AdvancedSceneManager.Editor.Popup<T>.overlay","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).overlay","nameWithType":"Popup<T>.overlay","nameWithType.vb":"Popup(Of T).overlay"},{"uid":"AdvancedSceneManager.Editor.Popup`1.rootVisualElement","name":"rootVisualElement","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_rootVisualElement","commentId":"F:AdvancedSceneManager.Editor.Popup`1.rootVisualElement","fullName":"AdvancedSceneManager.Editor.Popup<T>.rootVisualElement","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).rootVisualElement","nameWithType":"Popup<T>.rootVisualElement","nameWithType.vb":"Popup(Of T).rootVisualElement"},{"uid":"AdvancedSceneManager.Editor.Popup`1.isMainContentLoaded","name":"isMainContentLoaded","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_isMainContentLoaded","commentId":"P:AdvancedSceneManager.Editor.Popup`1.isMainContentLoaded","fullName":"AdvancedSceneManager.Editor.Popup<T>.isMainContentLoaded","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).isMainContentLoaded","nameWithType":"Popup<T>.isMainContentLoaded","nameWithType.vb":"Popup(Of T).isMainContentLoaded"},{"uid":"AdvancedSceneManager.Editor.Popup`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement)","name":"LoadContent(String, VisualElement)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_LoadContent_System_String_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.Popup<T>.LoadContent(System.String, UnityEngine.UIElements.VisualElement)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).LoadContent(System.String, UnityEngine.UIElements.VisualElement)","nameWithType":"Popup<T>.LoadContent(String, VisualElement)","nameWithType.vb":"Popup(Of T).LoadContent(String, VisualElement)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement,System.Boolean,System.Boolean,System.Boolean)","name":"LoadContent(String, VisualElement, Boolean, Boolean, Boolean)","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_LoadContent_System_String_UnityEngine_UIElements_VisualElement_System_Boolean_System_Boolean_System_Boolean_","commentId":"M:AdvancedSceneManager.Editor.Popup`1.LoadContent(System.String,UnityEngine.UIElements.VisualElement,System.Boolean,System.Boolean,System.Boolean)","fullName":"AdvancedSceneManager.Editor.Popup<T>.LoadContent(System.String, UnityEngine.UIElements.VisualElement, System.Boolean, System.Boolean, System.Boolean)","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).LoadContent(System.String, UnityEngine.UIElements.VisualElement, System.Boolean, System.Boolean, System.Boolean)","nameWithType":"Popup<T>.LoadContent(String, VisualElement, Boolean, Boolean, Boolean)","nameWithType.vb":"Popup(Of T).LoadContent(String, VisualElement, Boolean, Boolean, Boolean)"},{"uid":"AdvancedSceneManager.Editor.Popup`1.ReloadContent","name":"ReloadContent()","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_ReloadContent","commentId":"M:AdvancedSceneManager.Editor.Popup`1.ReloadContent","fullName":"AdvancedSceneManager.Editor.Popup<T>.ReloadContent()","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).ReloadContent()","nameWithType":"Popup<T>.ReloadContent()","nameWithType.vb":"Popup(Of T).ReloadContent()"},{"uid":"AdvancedSceneManager.Editor.Popup`1.enableBorder","name":"enableBorder","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_enableBorder","commentId":"P:AdvancedSceneManager.Editor.Popup`1.enableBorder","fullName":"AdvancedSceneManager.Editor.Popup<T>.enableBorder","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).enableBorder","nameWithType":"Popup<T>.enableBorder","nameWithType.vb":"Popup(Of T).enableBorder"},{"uid":"AdvancedSceneManager.Editor.Popup`1.hasBorder","name":"hasBorder","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_hasBorder","commentId":"P:AdvancedSceneManager.Editor.Popup`1.hasBorder","fullName":"AdvancedSceneManager.Editor.Popup<T>.hasBorder","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).hasBorder","nameWithType":"Popup<T>.hasBorder","nameWithType.vb":"Popup(Of T).hasBorder"},{"uid":"AdvancedSceneManager.Editor.Popup`1.offset","name":"offset","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_offset","commentId":"P:AdvancedSceneManager.Editor.Popup`1.offset","fullName":"AdvancedSceneManager.Editor.Popup<T>.offset","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).offset","nameWithType":"Popup<T>.offset","nameWithType.vb":"Popup(Of T).offset"},{"uid":"AdvancedSceneManager.Editor.Popup`1.alignRight","name":"alignRight","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_alignRight","commentId":"P:AdvancedSceneManager.Editor.Popup`1.alignRight","fullName":"AdvancedSceneManager.Editor.Popup<T>.alignRight","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).alignRight","nameWithType":"Popup<T>.alignRight","nameWithType.vb":"Popup(Of T).alignRight"},{"uid":"AdvancedSceneManager.Editor.Popup`1.placementTarget","name":"placementTarget","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_placementTarget","commentId":"P:AdvancedSceneManager.Editor.Popup`1.placementTarget","fullName":"AdvancedSceneManager.Editor.Popup<T>.placementTarget","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).placementTarget","nameWithType":"Popup<T>.placementTarget","nameWithType.vb":"Popup(Of T).placementTarget"},{"uid":"AdvancedSceneManager.Editor.Popup`1.parent","name":"parent","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_parent","commentId":"P:AdvancedSceneManager.Editor.Popup`1.parent","fullName":"AdvancedSceneManager.Editor.Popup<T>.parent","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).parent","nameWithType":"Popup<T>.parent","nameWithType.vb":"Popup(Of T).parent"},{"uid":"AdvancedSceneManager.Editor.Popup`1.SetPosition","name":"SetPosition()","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_SetPosition","commentId":"M:AdvancedSceneManager.Editor.Popup`1.SetPosition","fullName":"AdvancedSceneManager.Editor.Popup<T>.SetPosition()","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).SetPosition()","nameWithType":"Popup<T>.SetPosition()","nameWithType.vb":"Popup(Of T).SetPosition()"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Reopen*","name":"Reopen","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Reopen_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.Reopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.Reopen","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Reopen","nameWithType":"Popup<T>.Reopen","nameWithType.vb":"Popup(Of T).Reopen"},{"uid":"AdvancedSceneManager.Editor.Popup`1.OnReopen*","name":"OnReopen","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_OnReopen_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.OnReopen","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.OnReopen","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).OnReopen","nameWithType":"Popup<T>.OnReopen","nameWithType.vb":"Popup(Of T).OnReopen"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Open*","name":"Open","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Open_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.Open","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.Open","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Open","nameWithType":"Popup<T>.Open","nameWithType.vb":"Popup(Of T).Open"},{"uid":"AdvancedSceneManager.Editor.Popup`1.CloseWithoutAnimation*","name":"CloseWithoutAnimation","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_CloseWithoutAnimation_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.CloseWithoutAnimation","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.CloseWithoutAnimation","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).CloseWithoutAnimation","nameWithType":"Popup<T>.CloseWithoutAnimation","nameWithType.vb":"Popup(Of T).CloseWithoutAnimation"},{"uid":"AdvancedSceneManager.Editor.Popup`1.Close*","name":"Close","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_Close_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.Close","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.Close","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).Close","nameWithType":"Popup<T>.Close","nameWithType.vb":"Popup(Of T).Close"},{"uid":"AdvancedSceneManager.Editor.Popup`1.OnClose*","name":"OnClose","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_OnClose_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.OnClose","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.OnClose","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).OnClose","nameWithType":"Popup<T>.OnClose","nameWithType.vb":"Popup(Of T).OnClose"},{"uid":"AdvancedSceneManager.Editor.Popup`1.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_path_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.path","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).path","nameWithType":"Popup<T>.path","nameWithType.vb":"Popup(Of T).path"},{"uid":"AdvancedSceneManager.Editor.Popup`1.isMainContentLoaded*","name":"isMainContentLoaded","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_isMainContentLoaded_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.isMainContentLoaded","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.isMainContentLoaded","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).isMainContentLoaded","nameWithType":"Popup<T>.isMainContentLoaded","nameWithType.vb":"Popup(Of T).isMainContentLoaded"},{"uid":"AdvancedSceneManager.Editor.Popup`1.LoadContent*","name":"LoadContent","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_LoadContent_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.LoadContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.LoadContent","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).LoadContent","nameWithType":"Popup<T>.LoadContent","nameWithType.vb":"Popup(Of T).LoadContent"},{"uid":"AdvancedSceneManager.Editor.Popup`1.ReloadContent*","name":"ReloadContent","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_ReloadContent_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.ReloadContent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.ReloadContent","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).ReloadContent","nameWithType":"Popup<T>.ReloadContent","nameWithType.vb":"Popup(Of T).ReloadContent"},{"uid":"AdvancedSceneManager.Editor.Popup`1.enableBorder*","name":"enableBorder","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_enableBorder_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.enableBorder","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.enableBorder","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).enableBorder","nameWithType":"Popup<T>.enableBorder","nameWithType.vb":"Popup(Of T).enableBorder"},{"uid":"AdvancedSceneManager.Editor.Popup`1.hasBorder*","name":"hasBorder","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_hasBorder_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.hasBorder","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.hasBorder","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).hasBorder","nameWithType":"Popup<T>.hasBorder","nameWithType.vb":"Popup(Of T).hasBorder"},{"uid":"AdvancedSceneManager.Editor.Popup`1.offset*","name":"offset","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_offset_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.offset","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.offset","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).offset","nameWithType":"Popup<T>.offset","nameWithType.vb":"Popup(Of T).offset"},{"uid":"AdvancedSceneManager.Editor.Popup`1.alignRight*","name":"alignRight","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_alignRight_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.alignRight","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.alignRight","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).alignRight","nameWithType":"Popup<T>.alignRight","nameWithType.vb":"Popup(Of T).alignRight"},{"uid":"AdvancedSceneManager.Editor.Popup`1.placementTarget*","name":"placementTarget","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_placementTarget_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.placementTarget","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.placementTarget","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).placementTarget","nameWithType":"Popup<T>.placementTarget","nameWithType.vb":"Popup(Of T).placementTarget"},{"uid":"AdvancedSceneManager.Editor.Popup`1.parent*","name":"parent","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_parent_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.parent","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.parent","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).parent","nameWithType":"Popup<T>.parent","nameWithType.vb":"Popup(Of T).parent"},{"uid":"AdvancedSceneManager.Editor.Popup`1.SetPosition*","name":"SetPosition","href":"~/api/AdvancedSceneManager.Editor.Popup-1.yml#AdvancedSceneManager_Editor_Popup_1_SetPosition_","commentId":"Overload:AdvancedSceneManager.Editor.Popup`1.SetPosition","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Popup<T>.SetPosition","fullName.vb":"AdvancedSceneManager.Editor.Popup(Of T).SetPosition","nameWithType":"Popup<T>.SetPosition","nameWithType.vb":"Popup(Of T).SetPosition"}],"api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml":[{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlTraits","name":"SceneField.UxmlTraits","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml","commentId":"T:AdvancedSceneManager.Editor.SceneField.UxmlTraits","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlTraits","nameWithType":"SceneField.UxmlTraits"},{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription","name":"uxmlChildElementsDescription","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml#AdvancedSceneManager_Editor_SceneField_UxmlTraits_uxmlChildElementsDescription","commentId":"P:AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription","nameWithType":"SceneField.UxmlTraits.uxmlChildElementsDescription"},{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement,UnityEngine.UIElements.IUxmlAttributes,UnityEngine.UIElements.CreationContext)","name":"Init(VisualElement, IUxmlAttributes, CreationContext)","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml#AdvancedSceneManager_Editor_SceneField_UxmlTraits_Init_UnityEngine_UIElements_VisualElement_UnityEngine_UIElements_IUxmlAttributes_UnityEngine_UIElements_CreationContext_","commentId":"M:AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement,UnityEngine.UIElements.IUxmlAttributes,UnityEngine.UIElements.CreationContext)","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init(UnityEngine.UIElements.VisualElement, UnityEngine.UIElements.IUxmlAttributes, UnityEngine.UIElements.CreationContext)","nameWithType":"SceneField.UxmlTraits.Init(VisualElement, IUxmlAttributes, CreationContext)"},{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription*","name":"uxmlChildElementsDescription","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml#AdvancedSceneManager_Editor_SceneField_UxmlTraits_uxmlChildElementsDescription_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.uxmlChildElementsDescription","nameWithType":"SceneField.UxmlTraits.uxmlChildElementsDescription"},{"uid":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init*","name":"Init","href":"~/api/AdvancedSceneManager.Editor.SceneField.UxmlTraits.yml#AdvancedSceneManager_Editor_SceneField_UxmlTraits_Init_","commentId":"Overload:AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneField.UxmlTraits.Init","nameWithType":"SceneField.UxmlTraits.Init"}],"api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml":[{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow","name":"SceneOverviewWindow","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml","commentId":"T:AdvancedSceneManager.Editor.SceneOverviewWindow","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow","nameWithType":"SceneOverviewWindow"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.path","name":"path","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_path","commentId":"P:AdvancedSceneManager.Editor.SceneOverviewWindow.path","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.path","nameWithType":"SceneOverviewWindow.path"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_autoReloadOnWindowFocus","commentId":"P:AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus","nameWithType":"SceneOverviewWindow.autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable","name":"OnEnable()","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_OnEnable","commentId":"M:AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable()","nameWithType":"SceneOverviewWindow.OnEnable()"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.path*","name":"path","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_path_","commentId":"Overload:AdvancedSceneManager.Editor.SceneOverviewWindow.path","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.path","nameWithType":"SceneOverviewWindow.path"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus*","name":"autoReloadOnWindowFocus","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_autoReloadOnWindowFocus_","commentId":"Overload:AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.autoReloadOnWindowFocus","nameWithType":"SceneOverviewWindow.autoReloadOnWindowFocus"},{"uid":"AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.SceneOverviewWindow.yml#AdvancedSceneManager_Editor_SceneOverviewWindow_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.SceneOverviewWindow.OnEnable","nameWithType":"SceneOverviewWindow.OnEnable"}],"api/AdvancedSceneManager.Editor.TagsTab.yml":[{"uid":"AdvancedSceneManager.Editor.TagsTab","name":"TagsTab","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml","commentId":"T:AdvancedSceneManager.Editor.TagsTab","fullName":"AdvancedSceneManager.Editor.TagsTab","nameWithType":"TagsTab"},{"uid":"AdvancedSceneManager.Editor.TagsTab.OnEnable(UnityEngine.UIElements.VisualElement)","name":"OnEnable(VisualElement)","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_OnEnable_UnityEngine_UIElements_VisualElement_","commentId":"M:AdvancedSceneManager.Editor.TagsTab.OnEnable(UnityEngine.UIElements.VisualElement)","fullName":"AdvancedSceneManager.Editor.TagsTab.OnEnable(UnityEngine.UIElements.VisualElement)","nameWithType":"TagsTab.OnEnable(VisualElement)"},{"uid":"AdvancedSceneManager.Editor.TagsTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement,System.Int32)","name":"OnReorderEnd(SceneManagerWindow.DragAndDropReorder.DragElement, Int32)","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_OnReorderEnd_AdvancedSceneManager_Editor_SceneManagerWindow_DragAndDropReorder_DragElement_System_Int32_","commentId":"M:AdvancedSceneManager.Editor.TagsTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement,System.Int32)","fullName":"AdvancedSceneManager.Editor.TagsTab.OnReorderEnd(AdvancedSceneManager.Editor.SceneManagerWindow.DragAndDropReorder.DragElement, System.Int32)","nameWithType":"TagsTab.OnReorderEnd(SceneManagerWindow.DragAndDropReorder.DragElement, Int32)"},{"uid":"AdvancedSceneManager.Editor.TagsTab.FooterButtons","name":"FooterButtons","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_FooterButtons","commentId":"P:AdvancedSceneManager.Editor.TagsTab.FooterButtons","fullName":"AdvancedSceneManager.Editor.TagsTab.FooterButtons","nameWithType":"TagsTab.FooterButtons"},{"uid":"AdvancedSceneManager.Editor.TagsTab.OnEnable*","name":"OnEnable","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_OnEnable_","commentId":"Overload:AdvancedSceneManager.Editor.TagsTab.OnEnable","isSpec":"True","fullName":"AdvancedSceneManager.Editor.TagsTab.OnEnable","nameWithType":"TagsTab.OnEnable"},{"uid":"AdvancedSceneManager.Editor.TagsTab.OnReorderEnd*","name":"OnReorderEnd","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_OnReorderEnd_","commentId":"Overload:AdvancedSceneManager.Editor.TagsTab.OnReorderEnd","isSpec":"True","fullName":"AdvancedSceneManager.Editor.TagsTab.OnReorderEnd","nameWithType":"TagsTab.OnReorderEnd"},{"uid":"AdvancedSceneManager.Editor.TagsTab.FooterButtons*","name":"FooterButtons","href":"~/api/AdvancedSceneManager.Editor.TagsTab.yml#AdvancedSceneManager_Editor_TagsTab_FooterButtons_","commentId":"Overload:AdvancedSceneManager.Editor.TagsTab.FooterButtons","isSpec":"True","fullName":"AdvancedSceneManager.Editor.TagsTab.FooterButtons","nameWithType":"TagsTab.FooterButtons"}],"api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml":[{"uid":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility","name":"AssetDatabaseUtility","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml","commentId":"T:AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility","fullName":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility","nameWithType":"AssetDatabaseUtility"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh(System.Object)","name":"DisallowAutoRefresh(Object)","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml#AdvancedSceneManager_Editor_Utility_AssetDatabaseUtility_DisallowAutoRefresh_System_Object_","commentId":"M:AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh(System.Object)","fullName":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh(System.Object)","nameWithType":"AssetDatabaseUtility.DisallowAutoRefresh(Object)"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh(System.Object)","name":"AllowAutoRefresh(Object)","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml#AdvancedSceneManager_Editor_Utility_AssetDatabaseUtility_AllowAutoRefresh_System_Object_","commentId":"M:AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh(System.Object)","fullName":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh(System.Object)","nameWithType":"AssetDatabaseUtility.AllowAutoRefresh(Object)"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh*","name":"DisallowAutoRefresh","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml#AdvancedSceneManager_Editor_Utility_AssetDatabaseUtility_DisallowAutoRefresh_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.DisallowAutoRefresh","nameWithType":"AssetDatabaseUtility.DisallowAutoRefresh"},{"uid":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh*","name":"AllowAutoRefresh","href":"~/api/AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.yml#AdvancedSceneManager_Editor_Utility_AssetDatabaseUtility_AllowAutoRefresh_","commentId":"Overload:AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh","isSpec":"True","fullName":"AdvancedSceneManager.Editor.Utility.AssetDatabaseUtility.AllowAutoRefresh","nameWithType":"AssetDatabaseUtility.AllowAutoRefresh"}],"api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml":[{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy","name":"ASMSettings.SettingsProxy","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml","commentId":"T:AdvancedSceneManager.Models.ASMSettings.SettingsProxy","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy","nameWithType":"ASMSettings.SettingsProxy"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local","name":"local","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_local","commentId":"P:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local","nameWithType":"ASMSettings.SettingsProxy.local"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project","name":"project","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_project","commentId":"P:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project","nameWithType":"ASMSettings.SettingsProxy.project"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile","name":"profile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_profile","commentId":"P:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile","nameWithType":"ASMSettings.SettingsProxy.profile"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local*","name":"local","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_local_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.local","nameWithType":"ASMSettings.SettingsProxy.local"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project*","name":"project","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_project_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.project","nameWithType":"ASMSettings.SettingsProxy.project"},{"uid":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile*","name":"profile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.SettingsProxy.yml#AdvancedSceneManager_Models_ASMSettings_SettingsProxy_profile_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.SettingsProxy.profile","nameWithType":"ASMSettings.SettingsProxy.profile"}],"api/AdvancedSceneManager.Models.ASMSettings.yml":[{"uid":"AdvancedSceneManager.Models.ASMSettings","name":"ASMSettings","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml","commentId":"T:AdvancedSceneManager.Models.ASMSettings","fullName":"AdvancedSceneManager.Models.ASMSettings","nameWithType":"ASMSettings"},{"uid":"AdvancedSceneManager.Models.ASMSettings.profile","name":"profile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_profile","commentId":"P:AdvancedSceneManager.Models.ASMSettings.profile","fullName":"AdvancedSceneManager.Models.ASMSettings.profile","nameWithType":"ASMSettings.profile"},{"uid":"AdvancedSceneManager.Models.ASMSettings.buildProfile","name":"buildProfile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_buildProfile","commentId":"P:AdvancedSceneManager.Models.ASMSettings.buildProfile","fullName":"AdvancedSceneManager.Models.ASMSettings.buildProfile","nameWithType":"ASMSettings.buildProfile"},{"uid":"AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor","name":"buildUnitySplashScreenColor","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_buildUnitySplashScreenColor","commentId":"P:AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor","fullName":"AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor","nameWithType":"ASMSettings.buildUnitySplashScreenColor"},{"uid":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled","name":"inGameToolbarEnabled","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_inGameToolbarEnabled","commentId":"P:AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled","fullName":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled","nameWithType":"ASMSettings.inGameToolbarEnabled"},{"uid":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault","name":"inGameToolbarExpandedByDefault","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_inGameToolbarExpandedByDefault","commentId":"P:AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault","fullName":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault","nameWithType":"ASMSettings.inGameToolbarExpandedByDefault"},{"uid":"AdvancedSceneManager.Models.ASMSettings.name","name":"name","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_name","commentId":"P:AdvancedSceneManager.Models.ASMSettings.name","fullName":"AdvancedSceneManager.Models.ASMSettings.name","nameWithType":"ASMSettings.name"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Save","name":"Save()","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_Save","commentId":"M:AdvancedSceneManager.Models.ASMSettings.Save","fullName":"AdvancedSceneManager.Models.ASMSettings.Save()","nameWithType":"ASMSettings.Save()"},{"uid":"AdvancedSceneManager.Models.ASMSettings.MarkAsDirty","name":"MarkAsDirty()","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_MarkAsDirty","commentId":"M:AdvancedSceneManager.Models.ASMSettings.MarkAsDirty","fullName":"AdvancedSceneManager.Models.ASMSettings.MarkAsDirty()","nameWithType":"ASMSettings.MarkAsDirty()"},{"uid":"AdvancedSceneManager.Models.ASMSettings.profile*","name":"profile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_profile_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.profile","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.profile","nameWithType":"ASMSettings.profile"},{"uid":"AdvancedSceneManager.Models.ASMSettings.buildProfile*","name":"buildProfile","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_buildProfile_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.buildProfile","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.buildProfile","nameWithType":"ASMSettings.buildProfile"},{"uid":"AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor*","name":"buildUnitySplashScreenColor","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_buildUnitySplashScreenColor_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.buildUnitySplashScreenColor","nameWithType":"ASMSettings.buildUnitySplashScreenColor"},{"uid":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled*","name":"inGameToolbarEnabled","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_inGameToolbarEnabled_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarEnabled","nameWithType":"ASMSettings.inGameToolbarEnabled"},{"uid":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault*","name":"inGameToolbarExpandedByDefault","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_inGameToolbarExpandedByDefault_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.inGameToolbarExpandedByDefault","nameWithType":"ASMSettings.inGameToolbarExpandedByDefault"},{"uid":"AdvancedSceneManager.Models.ASMSettings.name*","name":"name","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_name_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.name","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.name","nameWithType":"ASMSettings.name"},{"uid":"AdvancedSceneManager.Models.ASMSettings.Save*","name":"Save","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_Save_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.Save","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.Save","nameWithType":"ASMSettings.Save"},{"uid":"AdvancedSceneManager.Models.ASMSettings.MarkAsDirty*","name":"MarkAsDirty","href":"~/api/AdvancedSceneManager.Models.ASMSettings.yml#AdvancedSceneManager_Models_ASMSettings_MarkAsDirty_","commentId":"Overload:AdvancedSceneManager.Models.ASMSettings.MarkAsDirty","isSpec":"True","fullName":"AdvancedSceneManager.Models.ASMSettings.MarkAsDirty","nameWithType":"ASMSettings.MarkAsDirty"}],"api/AdvancedSceneManager.Models.SceneTag.yml":[{"uid":"AdvancedSceneManager.Models.SceneTag","name":"SceneTag","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml","commentId":"T:AdvancedSceneManager.Models.SceneTag","fullName":"AdvancedSceneManager.Models.SceneTag","nameWithType":"SceneTag"},{"uid":"AdvancedSceneManager.Models.SceneTag.Default","name":"Default","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Default","commentId":"F:AdvancedSceneManager.Models.SceneTag.Default","fullName":"AdvancedSceneManager.Models.SceneTag.Default","nameWithType":"SceneTag.Default"},{"uid":"AdvancedSceneManager.Models.SceneTag.DoNotOpen","name":"DoNotOpen","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_DoNotOpen","commentId":"F:AdvancedSceneManager.Models.SceneTag.DoNotOpen","fullName":"AdvancedSceneManager.Models.SceneTag.DoNotOpen","nameWithType":"SceneTag.DoNotOpen"},{"uid":"AdvancedSceneManager.Models.SceneTag.Persistent","name":"Persistent","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Persistent","commentId":"F:AdvancedSceneManager.Models.SceneTag.Persistent","fullName":"AdvancedSceneManager.Models.SceneTag.Persistent","nameWithType":"SceneTag.Persistent"},{"uid":"AdvancedSceneManager.Models.SceneTag.PersistIfRequired","name":"PersistIfRequired","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_PersistIfRequired","commentId":"F:AdvancedSceneManager.Models.SceneTag.PersistIfRequired","fullName":"AdvancedSceneManager.Models.SceneTag.PersistIfRequired","nameWithType":"SceneTag.PersistIfRequired"},{"uid":"AdvancedSceneManager.Models.SceneTag.#ctor","name":"SceneTag()","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag__ctor","commentId":"M:AdvancedSceneManager.Models.SceneTag.#ctor","fullName":"AdvancedSceneManager.Models.SceneTag.SceneTag()","nameWithType":"SceneTag.SceneTag()"},{"uid":"AdvancedSceneManager.Models.SceneTag.#ctor(System.String,System.Nullable{UnityEngine.Color},System.String)","name":"SceneTag(String, Nullable<Color>, String)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag__ctor_System_String_System_Nullable_UnityEngine_Color__System_String_","commentId":"M:AdvancedSceneManager.Models.SceneTag.#ctor(System.String,System.Nullable{UnityEngine.Color},System.String)","name.vb":"SceneTag(String, Nullable(Of Color), String)","fullName":"AdvancedSceneManager.Models.SceneTag.SceneTag(System.String, System.Nullable<UnityEngine.Color>, System.String)","fullName.vb":"AdvancedSceneManager.Models.SceneTag.SceneTag(System.String, System.Nullable(Of UnityEngine.Color), System.String)","nameWithType":"SceneTag.SceneTag(String, Nullable<Color>, String)","nameWithType.vb":"SceneTag.SceneTag(String, Nullable(Of Color), String)"},{"uid":"AdvancedSceneManager.Models.SceneTag.name","name":"name","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_name","commentId":"F:AdvancedSceneManager.Models.SceneTag.name","fullName":"AdvancedSceneManager.Models.SceneTag.name","nameWithType":"SceneTag.name"},{"uid":"AdvancedSceneManager.Models.SceneTag.label","name":"label","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_label","commentId":"F:AdvancedSceneManager.Models.SceneTag.label","fullName":"AdvancedSceneManager.Models.SceneTag.label","nameWithType":"SceneTag.label"},{"uid":"AdvancedSceneManager.Models.SceneTag.id","name":"id","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_id","commentId":"F:AdvancedSceneManager.Models.SceneTag.id","fullName":"AdvancedSceneManager.Models.SceneTag.id","nameWithType":"SceneTag.id"},{"uid":"AdvancedSceneManager.Models.SceneTag.color","name":"color","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_color","commentId":"F:AdvancedSceneManager.Models.SceneTag.color","fullName":"AdvancedSceneManager.Models.SceneTag.color","nameWithType":"SceneTag.color"},{"uid":"AdvancedSceneManager.Models.SceneTag.closeBehavior","name":"closeBehavior","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_closeBehavior","commentId":"F:AdvancedSceneManager.Models.SceneTag.closeBehavior","fullName":"AdvancedSceneManager.Models.SceneTag.closeBehavior","nameWithType":"SceneTag.closeBehavior"},{"uid":"AdvancedSceneManager.Models.SceneTag.openBehavior","name":"openBehavior","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_openBehavior","commentId":"F:AdvancedSceneManager.Models.SceneTag.openBehavior","fullName":"AdvancedSceneManager.Models.SceneTag.openBehavior","nameWithType":"SceneTag.openBehavior"},{"uid":"AdvancedSceneManager.Models.SceneTag.Find(System.String)","name":"Find(String)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Find_System_String_","commentId":"M:AdvancedSceneManager.Models.SceneTag.Find(System.String)","fullName":"AdvancedSceneManager.Models.SceneTag.Find(System.String)","nameWithType":"SceneTag.Find(String)"},{"uid":"AdvancedSceneManager.Models.SceneTag.Equals(System.Object)","name":"Equals(Object)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Equals_System_Object_","commentId":"M:AdvancedSceneManager.Models.SceneTag.Equals(System.Object)","fullName":"AdvancedSceneManager.Models.SceneTag.Equals(System.Object)","nameWithType":"SceneTag.Equals(Object)"},{"uid":"AdvancedSceneManager.Models.SceneTag.GetHashCode","name":"GetHashCode()","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_GetHashCode","commentId":"M:AdvancedSceneManager.Models.SceneTag.GetHashCode","fullName":"AdvancedSceneManager.Models.SceneTag.GetHashCode()","nameWithType":"SceneTag.GetHashCode()"},{"uid":"AdvancedSceneManager.Models.SceneTag.Equals(AdvancedSceneManager.Models.SceneTag)","name":"Equals(SceneTag)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Equals_AdvancedSceneManager_Models_SceneTag_","commentId":"M:AdvancedSceneManager.Models.SceneTag.Equals(AdvancedSceneManager.Models.SceneTag)","fullName":"AdvancedSceneManager.Models.SceneTag.Equals(AdvancedSceneManager.Models.SceneTag)","nameWithType":"SceneTag.Equals(SceneTag)"},{"uid":"AdvancedSceneManager.Models.SceneTag.op_Equality(AdvancedSceneManager.Models.SceneTag,AdvancedSceneManager.Models.SceneTag)","name":"Equality(SceneTag, SceneTag)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_op_Equality_AdvancedSceneManager_Models_SceneTag_AdvancedSceneManager_Models_SceneTag_","commentId":"M:AdvancedSceneManager.Models.SceneTag.op_Equality(AdvancedSceneManager.Models.SceneTag,AdvancedSceneManager.Models.SceneTag)","fullName":"AdvancedSceneManager.Models.SceneTag.Equality(AdvancedSceneManager.Models.SceneTag, AdvancedSceneManager.Models.SceneTag)","nameWithType":"SceneTag.Equality(SceneTag, SceneTag)"},{"uid":"AdvancedSceneManager.Models.SceneTag.op_Inequality(AdvancedSceneManager.Models.SceneTag,AdvancedSceneManager.Models.SceneTag)","name":"Inequality(SceneTag, SceneTag)","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_op_Inequality_AdvancedSceneManager_Models_SceneTag_AdvancedSceneManager_Models_SceneTag_","commentId":"M:AdvancedSceneManager.Models.SceneTag.op_Inequality(AdvancedSceneManager.Models.SceneTag,AdvancedSceneManager.Models.SceneTag)","fullName":"AdvancedSceneManager.Models.SceneTag.Inequality(AdvancedSceneManager.Models.SceneTag, AdvancedSceneManager.Models.SceneTag)","nameWithType":"SceneTag.Inequality(SceneTag, SceneTag)"},{"uid":"AdvancedSceneManager.Models.SceneTag.ToString","name":"ToString()","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_ToString","commentId":"M:AdvancedSceneManager.Models.SceneTag.ToString","fullName":"AdvancedSceneManager.Models.SceneTag.ToString()","nameWithType":"SceneTag.ToString()"},{"uid":"AdvancedSceneManager.Models.SceneTag.#ctor*","name":"SceneTag","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag__ctor_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.#ctor","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.SceneTag","nameWithType":"SceneTag.SceneTag"},{"uid":"AdvancedSceneManager.Models.SceneTag.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Find_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.Find","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.Find","nameWithType":"SceneTag.Find"},{"uid":"AdvancedSceneManager.Models.SceneTag.Equals*","name":"Equals","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_Equals_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.Equals","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.Equals","nameWithType":"SceneTag.Equals"},{"uid":"AdvancedSceneManager.Models.SceneTag.GetHashCode*","name":"GetHashCode","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_GetHashCode_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.GetHashCode","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.GetHashCode","nameWithType":"SceneTag.GetHashCode"},{"uid":"AdvancedSceneManager.Models.SceneTag.op_Equality*","name":"Equality","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_op_Equality_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.op_Equality","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.Equality","nameWithType":"SceneTag.Equality"},{"uid":"AdvancedSceneManager.Models.SceneTag.op_Inequality*","name":"Inequality","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_op_Inequality_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.op_Inequality","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.Inequality","nameWithType":"SceneTag.Inequality"},{"uid":"AdvancedSceneManager.Models.SceneTag.ToString*","name":"ToString","href":"~/api/AdvancedSceneManager.Models.SceneTag.yml#AdvancedSceneManager_Models_SceneTag_ToString_","commentId":"Overload:AdvancedSceneManager.Models.SceneTag.ToString","isSpec":"True","fullName":"AdvancedSceneManager.Models.SceneTag.ToString","nameWithType":"SceneTag.ToString"}],"api/AdvancedSceneManager.Models.TagList.yml":[{"uid":"AdvancedSceneManager.Models.TagList","name":"TagList","href":"~/api/AdvancedSceneManager.Models.TagList.yml","commentId":"T:AdvancedSceneManager.Models.TagList","fullName":"AdvancedSceneManager.Models.TagList","nameWithType":"TagList"},{"uid":"AdvancedSceneManager.Models.TagList.Item(System.String)","name":"Item[String]","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_Item_System_String_","commentId":"P:AdvancedSceneManager.Models.TagList.Item(System.String)","name.vb":"Item(String)","fullName":"AdvancedSceneManager.Models.TagList.Item[System.String]","fullName.vb":"AdvancedSceneManager.Models.TagList.Item(System.String)","nameWithType":"TagList.Item[String]","nameWithType.vb":"TagList.Item(String)"},{"uid":"AdvancedSceneManager.Models.TagList.Item(AdvancedSceneManager.Models.Scene)","name":"Item[Scene]","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_Item_AdvancedSceneManager_Models_Scene_","commentId":"P:AdvancedSceneManager.Models.TagList.Item(AdvancedSceneManager.Models.Scene)","name.vb":"Item(Scene)","fullName":"AdvancedSceneManager.Models.TagList.Item[AdvancedSceneManager.Models.Scene]","fullName.vb":"AdvancedSceneManager.Models.TagList.Item(AdvancedSceneManager.Models.Scene)","nameWithType":"TagList.Item[Scene]","nameWithType.vb":"TagList.Item(Scene)"},{"uid":"AdvancedSceneManager.Models.TagList.TryGetValue(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneTag@)","name":"TryGetValue(Scene, out SceneTag)","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_TryGetValue_AdvancedSceneManager_Models_Scene_AdvancedSceneManager_Models_SceneTag__","commentId":"M:AdvancedSceneManager.Models.TagList.TryGetValue(AdvancedSceneManager.Models.Scene,AdvancedSceneManager.Models.SceneTag@)","name.vb":"TryGetValue(Scene, ByRef SceneTag)","fullName":"AdvancedSceneManager.Models.TagList.TryGetValue(AdvancedSceneManager.Models.Scene, out AdvancedSceneManager.Models.SceneTag)","fullName.vb":"AdvancedSceneManager.Models.TagList.TryGetValue(AdvancedSceneManager.Models.Scene, ByRef AdvancedSceneManager.Models.SceneTag)","nameWithType":"TagList.TryGetValue(Scene, out SceneTag)","nameWithType.vb":"TagList.TryGetValue(Scene, ByRef SceneTag)"},{"uid":"AdvancedSceneManager.Models.TagList.TryGetValue(System.String,AdvancedSceneManager.Models.SceneTag@)","name":"TryGetValue(String, out SceneTag)","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_TryGetValue_System_String_AdvancedSceneManager_Models_SceneTag__","commentId":"M:AdvancedSceneManager.Models.TagList.TryGetValue(System.String,AdvancedSceneManager.Models.SceneTag@)","name.vb":"TryGetValue(String, ByRef SceneTag)","fullName":"AdvancedSceneManager.Models.TagList.TryGetValue(System.String, out AdvancedSceneManager.Models.SceneTag)","fullName.vb":"AdvancedSceneManager.Models.TagList.TryGetValue(System.String, ByRef AdvancedSceneManager.Models.SceneTag)","nameWithType":"TagList.TryGetValue(String, out SceneTag)","nameWithType.vb":"TagList.TryGetValue(String, ByRef SceneTag)"},{"uid":"AdvancedSceneManager.Models.TagList.Item*","name":"Item","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_Item_","commentId":"Overload:AdvancedSceneManager.Models.TagList.Item","isSpec":"True","fullName":"AdvancedSceneManager.Models.TagList.Item","nameWithType":"TagList.Item"},{"uid":"AdvancedSceneManager.Models.TagList.TryGetValue*","name":"TryGetValue","href":"~/api/AdvancedSceneManager.Models.TagList.yml#AdvancedSceneManager_Models_TagList_TryGetValue_","commentId":"Overload:AdvancedSceneManager.Models.TagList.TryGetValue","isSpec":"True","fullName":"AdvancedSceneManager.Models.TagList.TryGetValue","nameWithType":"TagList.TryGetValue"}],"api/AdvancedSceneManager.Utility.GuidReference.yml":[{"uid":"AdvancedSceneManager.Utility.GuidReference","name":"GuidReference","href":"~/api/AdvancedSceneManager.Utility.GuidReference.yml","commentId":"T:AdvancedSceneManager.Utility.GuidReference","fullName":"AdvancedSceneManager.Utility.GuidReference","nameWithType":"GuidReference"},{"uid":"AdvancedSceneManager.Utility.GuidReference.guid","name":"guid","href":"~/api/AdvancedSceneManager.Utility.GuidReference.yml#AdvancedSceneManager_Utility_GuidReference_guid","commentId":"F:AdvancedSceneManager.Utility.GuidReference.guid","fullName":"AdvancedSceneManager.Utility.GuidReference.guid","nameWithType":"GuidReference.guid"}],"api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml":[{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility","name":"GuidReferenceUtility","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml","commentId":"T:AdvancedSceneManager.Utility.GuidReferenceUtility","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility","nameWithType":"GuidReferenceUtility"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime(UnityEngine.Object)","name":"AddRuntime(Object)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_AddRuntime_UnityEngine_Object_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime(UnityEngine.Object)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime(UnityEngine.Object)","nameWithType":"GuidReferenceUtility.AddRuntime(Object)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(UnityEngine.Object)","name":"RemoveRuntime(Object)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_RemoveRuntime_UnityEngine_Object_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(UnityEngine.Object)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(UnityEngine.Object)","nameWithType":"GuidReferenceUtility.RemoveRuntime(Object)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(System.String)","name":"RemoveRuntime(String)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_RemoveRuntime_System_String_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(System.String)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime(System.String)","nameWithType":"GuidReferenceUtility.RemoveRuntime(String)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference(System.String)","name":"HasReference(String)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_HasReference_System_String_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference(System.String)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference(System.String)","nameWithType":"GuidReferenceUtility.HasReference(String)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind``1(System.String,``0@)","name":"TryFind<T>(String, out T)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_TryFind__1_System_String___0__","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind``1(System.String,``0@)","name.vb":"TryFind(Of T)(String, ByRef T)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind<T>(System.String, out T)","fullName.vb":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind(Of T)(System.String, ByRef T)","nameWithType":"GuidReferenceUtility.TryFind<T>(String, out T)","nameWithType.vb":"GuidReferenceUtility.TryFind(Of T)(String, ByRef T)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind(System.String,UnityEngine.Object@)","name":"TryFind(String, out Object)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_TryFind_System_String_UnityEngine_Object__","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind(System.String,UnityEngine.Object@)","name.vb":"TryFind(String, ByRef Object)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind(System.String, out UnityEngine.Object)","fullName.vb":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind(System.String, ByRef UnityEngine.Object)","nameWithType":"GuidReferenceUtility.TryFind(String, out Object)","nameWithType.vb":"GuidReferenceUtility.TryFind(String, ByRef Object)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String)","name":"Find(String)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_Find_System_String_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String)","nameWithType":"GuidReferenceUtility.Find(String)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find``1(System.String)","name":"Find<T>(String)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_Find__1_System_String_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.Find``1(System.String)","name.vb":"Find(Of T)(String)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find<T>(System.String)","fullName.vb":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(Of T)(System.String)","nameWithType":"GuidReferenceUtility.Find<T>(String)","nameWithType.vb":"GuidReferenceUtility.Find(Of T)(String)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String,System.Action{UnityEngine.Object})","name":"Find(String, Action<Object>)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_Find_System_String_System_Action_UnityEngine_Object__","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String,System.Action{UnityEngine.Object})","name.vb":"Find(String, Action(Of Object))","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String, System.Action<UnityEngine.Object>)","fullName.vb":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find(System.String, System.Action(Of UnityEngine.Object))","nameWithType":"GuidReferenceUtility.Find(String, Action<Object>)","nameWithType.vb":"GuidReferenceUtility.Find(String, Action(Of Object))"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent(UnityEngine.GameObject)","name":"GetOrAddPersistent(GameObject)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_GetOrAddPersistent_UnityEngine_GameObject_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent(UnityEngine.GameObject)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent(UnityEngine.GameObject)","nameWithType":"GuidReferenceUtility.GetOrAddPersistent(GameObject)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent(UnityEngine.GameObject)","name":"AddPersistent(GameObject)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_AddPersistent_UnityEngine_GameObject_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent(UnityEngine.GameObject)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent(UnityEngine.GameObject)","nameWithType":"GuidReferenceUtility.AddPersistent(GameObject)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent(UnityEngine.GameObject,System.Boolean)","name":"RemovePersistent(GameObject, Boolean)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_RemovePersistent_UnityEngine_GameObject_System_Boolean_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent(UnityEngine.GameObject,System.Boolean)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent(UnityEngine.GameObject, System.Boolean)","nameWithType":"GuidReferenceUtility.RemovePersistent(GameObject, Boolean)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID","name":"GenerateID()","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_GenerateID","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID()","nameWithType":"GuidReferenceUtility.GenerateID()"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent(System.String)","name":"FindPersistent(String)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_FindPersistent_System_String_","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent(System.String)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent(System.String)","nameWithType":"GuidReferenceUtility.FindPersistent(String)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent(System.String,UnityEngine.GameObject@)","name":"TryFindPersistent(String, out GameObject)","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_TryFindPersistent_System_String_UnityEngine_GameObject__","commentId":"M:AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent(System.String,UnityEngine.GameObject@)","name.vb":"TryFindPersistent(String, ByRef GameObject)","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent(System.String, out UnityEngine.GameObject)","fullName.vb":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent(System.String, ByRef UnityEngine.GameObject)","nameWithType":"GuidReferenceUtility.TryFindPersistent(String, out GameObject)","nameWithType.vb":"GuidReferenceUtility.TryFindPersistent(String, ByRef GameObject)"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime*","name":"AddRuntime","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_AddRuntime_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddRuntime","nameWithType":"GuidReferenceUtility.AddRuntime"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime*","name":"RemoveRuntime","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_RemoveRuntime_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemoveRuntime","nameWithType":"GuidReferenceUtility.RemoveRuntime"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference*","name":"HasReference","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_HasReference_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.HasReference","nameWithType":"GuidReferenceUtility.HasReference"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind*","name":"TryFind","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_TryFind_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFind","nameWithType":"GuidReferenceUtility.TryFind"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find*","name":"Find","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_Find_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.Find","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.Find","nameWithType":"GuidReferenceUtility.Find"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent*","name":"GetOrAddPersistent","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_GetOrAddPersistent_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.GetOrAddPersistent","nameWithType":"GuidReferenceUtility.GetOrAddPersistent"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent*","name":"AddPersistent","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_AddPersistent_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.AddPersistent","nameWithType":"GuidReferenceUtility.AddPersistent"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent*","name":"RemovePersistent","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_RemovePersistent_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.RemovePersistent","nameWithType":"GuidReferenceUtility.RemovePersistent"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID*","name":"GenerateID","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_GenerateID_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.GenerateID","nameWithType":"GuidReferenceUtility.GenerateID"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent*","name":"FindPersistent","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_FindPersistent_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.FindPersistent","nameWithType":"GuidReferenceUtility.FindPersistent"},{"uid":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent*","name":"TryFindPersistent","href":"~/api/AdvancedSceneManager.Utility.GuidReferenceUtility.yml#AdvancedSceneManager_Utility_GuidReferenceUtility_TryFindPersistent_","commentId":"Overload:AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent","isSpec":"True","fullName":"AdvancedSceneManager.Utility.GuidReferenceUtility.TryFindPersistent","nameWithType":"GuidReferenceUtility.TryFindPersistent"}],"api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml":[{"uid":"AdvancedSceneManager.Utility.ScriptableObjectUtility","name":"ScriptableObjectUtility","href":"~/api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml","commentId":"T:AdvancedSceneManager.Utility.ScriptableObjectUtility","fullName":"AdvancedSceneManager.Utility.ScriptableObjectUtility","nameWithType":"ScriptableObjectUtility"},{"uid":"AdvancedSceneManager.Utility.ScriptableObjectUtility.Save(UnityEngine.ScriptableObject)","name":"Save(ScriptableObject)","href":"~/api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml#AdvancedSceneManager_Utility_ScriptableObjectUtility_Save_UnityEngine_ScriptableObject_","commentId":"M:AdvancedSceneManager.Utility.ScriptableObjectUtility.Save(UnityEngine.ScriptableObject)","fullName":"AdvancedSceneManager.Utility.ScriptableObjectUtility.Save(UnityEngine.ScriptableObject)","nameWithType":"ScriptableObjectUtility.Save(ScriptableObject)"},{"uid":"AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton``1(System.String,System.String)","name":"GetSingleton<T>(String, String)","href":"~/api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml#AdvancedSceneManager_Utility_ScriptableObjectUtility_GetSingleton__1_System_String_System_String_","commentId":"M:AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton``1(System.String,System.String)","name.vb":"GetSingleton(Of T)(String, String)","fullName":"AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton<T>(System.String, System.String)","fullName.vb":"AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton(Of T)(System.String, System.String)","nameWithType":"ScriptableObjectUtility.GetSingleton<T>(String, String)","nameWithType.vb":"ScriptableObjectUtility.GetSingleton(Of T)(String, String)"},{"uid":"AdvancedSceneManager.Utility.ScriptableObjectUtility.Save*","name":"Save","href":"~/api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml#AdvancedSceneManager_Utility_ScriptableObjectUtility_Save_","commentId":"Overload:AdvancedSceneManager.Utility.ScriptableObjectUtility.Save","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ScriptableObjectUtility.Save","nameWithType":"ScriptableObjectUtility.Save"},{"uid":"AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton*","name":"GetSingleton","href":"~/api/AdvancedSceneManager.Utility.ScriptableObjectUtility.yml#AdvancedSceneManager_Utility_ScriptableObjectUtility_GetSingleton_","commentId":"Overload:AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton","isSpec":"True","fullName":"AdvancedSceneManager.Utility.ScriptableObjectUtility.GetSingleton","nameWithType":"ScriptableObjectUtility.GetSingleton"}],"api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml":[{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2","name":"SerializableDictionary<TKey, TValue>","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml","commentId":"T:AdvancedSceneManager.Utility.SerializableDictionary`2","name.vb":"SerializableDictionary(Of TKey, TValue)","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue)","nameWithType":"SerializableDictionary<TKey, TValue>","nameWithType.vb":"SerializableDictionary(Of TKey, TValue)"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.throwOnDeserializeWhenKeyValueMismatch","name":"throwOnDeserializeWhenKeyValueMismatch","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_throwOnDeserializeWhenKeyValueMismatch","commentId":"P:AdvancedSceneManager.Utility.SerializableDictionary`2.throwOnDeserializeWhenKeyValueMismatch","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.throwOnDeserializeWhenKeyValueMismatch","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).throwOnDeserializeWhenKeyValueMismatch","nameWithType":"SerializableDictionary<TKey, TValue>.throwOnDeserializeWhenKeyValueMismatch","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).throwOnDeserializeWhenKeyValueMismatch"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.keys","name":"keys","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_keys","commentId":"F:AdvancedSceneManager.Utility.SerializableDictionary`2.keys","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.keys","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).keys","nameWithType":"SerializableDictionary<TKey, TValue>.keys","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).keys"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.values","name":"values","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_values","commentId":"F:AdvancedSceneManager.Utility.SerializableDictionary`2.values","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.values","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).values","nameWithType":"SerializableDictionary<TKey, TValue>.values","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).values"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.OnBeforeSerialize","name":"OnBeforeSerialize()","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_OnBeforeSerialize","commentId":"M:AdvancedSceneManager.Utility.SerializableDictionary`2.OnBeforeSerialize","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.OnBeforeSerialize()","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).OnBeforeSerialize()","nameWithType":"SerializableDictionary<TKey, TValue>.OnBeforeSerialize()","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).OnBeforeSerialize()"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.OnAfterDeserialize","name":"OnAfterDeserialize()","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_OnAfterDeserialize","commentId":"M:AdvancedSceneManager.Utility.SerializableDictionary`2.OnAfterDeserialize","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.OnAfterDeserialize()","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).OnAfterDeserialize()","nameWithType":"SerializableDictionary<TKey, TValue>.OnAfterDeserialize()","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).OnAfterDeserialize()"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.throwOnDeserializeWhenKeyValueMismatch*","name":"throwOnDeserializeWhenKeyValueMismatch","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_throwOnDeserializeWhenKeyValueMismatch_","commentId":"Overload:AdvancedSceneManager.Utility.SerializableDictionary`2.throwOnDeserializeWhenKeyValueMismatch","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.throwOnDeserializeWhenKeyValueMismatch","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).throwOnDeserializeWhenKeyValueMismatch","nameWithType":"SerializableDictionary<TKey, TValue>.throwOnDeserializeWhenKeyValueMismatch","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).throwOnDeserializeWhenKeyValueMismatch"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.OnBeforeSerialize*","name":"OnBeforeSerialize","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_OnBeforeSerialize_","commentId":"Overload:AdvancedSceneManager.Utility.SerializableDictionary`2.OnBeforeSerialize","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.OnBeforeSerialize","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).OnBeforeSerialize","nameWithType":"SerializableDictionary<TKey, TValue>.OnBeforeSerialize","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).OnBeforeSerialize"},{"uid":"AdvancedSceneManager.Utility.SerializableDictionary`2.OnAfterDeserialize*","name":"OnAfterDeserialize","href":"~/api/AdvancedSceneManager.Utility.SerializableDictionary-2.yml#AdvancedSceneManager_Utility_SerializableDictionary_2_OnAfterDeserialize_","commentId":"Overload:AdvancedSceneManager.Utility.SerializableDictionary`2.OnAfterDeserialize","isSpec":"True","fullName":"AdvancedSceneManager.Utility.SerializableDictionary<TKey, TValue>.OnAfterDeserialize","fullName.vb":"AdvancedSceneManager.Utility.SerializableDictionary(Of TKey, TValue).OnAfterDeserialize","nameWithType":"SerializableDictionary<TKey, TValue>.OnAfterDeserialize","nameWithType.vb":"SerializableDictionary(Of TKey, TValue).OnAfterDeserialize"}],"index.md":[],"guides/Profile.md":[],"guides/QuickStart.md":[],"guides/Callbacks.md":[],"guides/InGameToolbar.md":[],"guides/LoadingScreen.md":[],"guides/PauseScreenUtility.md":[],"guides/PreloadedSceneHelper.md":[],"guides/readme.md":[],"guides/Scene.md":[],"guides/SceneAction.md":[],"guides/SceneCollection.md":[],"guides/SceneHelper.md":[],"guides/SceneManager.md":[],"guides/SceneManagerWindow.md":[],"guides/SceneOperation.md":[],"guides/SceneOverviewWindow.md":[],"guides/SplashScreen.md":[],"plugins/plugin.asm.addressables.md":[],"plugins/plugin.asm.cross-scene-references.md":[],"plugins/plugin.asm.locking.md":[],"guides/toc.yml":[],"plugins/toc.yml":[],"toc.yml":[],"api/toc.yml":[],"image/merge-scenes-menu.png":[],"image/menu.png":[],"image/locking-warning.png":[],"image/in-game-toolbar.png":[],"image/quick-start-setup.png":[],"image/profile-dropdown.png":[],"image/package-manager.png":[],"image/package-manager-menu.png":[],"image/loading-screen-variables.png":[],"image/loading-screen-override.png":[],"image/guid-reference.png":[],"image/git-package-menu.png":[],"image/cross-scene-indicator.png":[],"image/cross-scene-debugger-menu.png":[],"image/coroutine-runner.png":[],"image/combine-scenes.png":[],"image/callback-analyzer-menu.png":[],"image/button-quit.png":[],"image/blacklist.png":[],"image/addressables.png":[],"image/=.png":[],"image/Unity-event.png":[],"image/tags.png":[],"image/split-scene-result.png":[],"image/settings.png":[],"image/settings-splashscreen.png":[],"image/selection.png":[],"image/scripting define symbols.png":[],"image/preload-example.png":[],"image/header.png":[],"resources/logo.png":[],"resources/icon.png":[],"resources/favicon.ico":[],"image/Scene-reference.png":[],"image/scene-overview.png":[],"image/scene-manager-menu.png":[],"image/scene-helper.png":[],"image/File-menu-and-scene-manager-window.png":[],"image/experimental-packages.png":[],"image/dynamic-collections.png":[],"image/cross-scene-reference.png":[],"image/cross-scene-reference-debugger2.png":[],"image/cross-scene-reference-debugger.png":[],"image/combine-scenes-result.png":[],"image/collection.png":[],"image/collection-edit-menu.png":[],"image/callbackutility.png":[],"image/button-open-collection.png":[],"image/bake-lightmaps.png":[],"image/+.png":[],"image/▶.png":[],"image/plugins-and-samples.PNG":[],"image/play.png":[],"image/pause-screen.png":[],"image/new-collection.png":[],"resources/ExampleScriptingApi.png":[],"resources/ExampleManual.png":[],"image/scenes.png":[],"image/scene-split-menu.png":[],"image/open.png":[],"image/new-tag.png":[],"image/locking-scene.png":[],"image/locking-collection.png":[],"image/-.png":[],"faq.md":[]}